VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram6t512x192
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 260.224 BY 105.792 ;
  SYMMETRY X Y R90 ;

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 237.120 0.000 237.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 237.120 0.000 237.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 237.120 0.000 237.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 237.120 0.000 237.272 0.152 ;
    END
  END CE1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 235.904 0.000 236.056 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 235.904 0.000 236.056 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 235.904 0.000 236.056 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 235.904 0.000 236.056 0.152 ;
    END
  END CSB1

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 234.688 0.000 234.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 234.688 0.000 234.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 234.688 0.000 234.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 234.688 0.000 234.840 0.152 ;
    END
  END OEB1

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 233.472 0.000 233.624 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 233.472 0.000 233.624 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 233.472 0.000 233.624 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 233.472 0.000 233.624 0.152 ;
    END
  END O1[3]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 233.168 0.000 233.320 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 233.168 0.000 233.320 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 233.168 0.000 233.320 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 233.168 0.000 233.320 0.152 ;
    END
  END O1[2]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 232.864 0.000 233.016 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 232.864 0.000 233.016 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 232.864 0.000 233.016 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 232.864 0.000 233.016 0.152 ;
    END
  END O1[1]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 232.560 0.000 232.712 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 232.560 0.000 232.712 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 232.560 0.000 232.712 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 232.560 0.000 232.712 0.152 ;
    END
  END O1[0]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 231.344 0.000 231.496 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 231.344 0.000 231.496 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 231.344 0.000 231.496 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 231.344 0.000 231.496 0.152 ;
    END
  END I1[0]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 231.040 0.000 231.192 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 231.040 0.000 231.192 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 231.040 0.000 231.192 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 231.040 0.000 231.192 0.152 ;
    END
  END I1[1]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 230.736 0.000 230.888 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 230.736 0.000 230.888 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 230.736 0.000 230.888 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 230.736 0.000 230.888 0.152 ;
    END
  END I1[2]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 230.432 0.000 230.584 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 230.432 0.000 230.584 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 230.432 0.000 230.584 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 230.432 0.000 230.584 0.152 ;
    END
  END I1[3]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 229.216 0.000 229.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 229.216 0.000 229.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 229.216 0.000 229.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 229.216 0.000 229.368 0.152 ;
    END
  END O1[7]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 228.912 0.000 229.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 228.912 0.000 229.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 228.912 0.000 229.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 228.912 0.000 229.064 0.152 ;
    END
  END O1[6]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 228.608 0.000 228.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 228.608 0.000 228.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 228.608 0.000 228.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 228.608 0.000 228.760 0.152 ;
    END
  END O1[5]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 228.304 0.000 228.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 228.304 0.000 228.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 228.304 0.000 228.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 228.304 0.000 228.456 0.152 ;
    END
  END O1[4]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 227.088 0.000 227.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 227.088 0.000 227.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 227.088 0.000 227.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 227.088 0.000 227.240 0.152 ;
    END
  END I1[4]

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.784 0.000 226.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 226.784 0.000 226.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 226.784 0.000 226.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 226.784 0.000 226.936 0.152 ;
    END
  END I1[5]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.480 0.000 226.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 226.480 0.000 226.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 226.480 0.000 226.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 226.480 0.000 226.632 0.152 ;
    END
  END I1[6]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.176 0.000 226.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 226.176 0.000 226.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 226.176 0.000 226.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 226.176 0.000 226.328 0.152 ;
    END
  END I1[7]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 224.960 0.000 225.112 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 224.960 0.000 225.112 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 224.960 0.000 225.112 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 224.960 0.000 225.112 0.152 ;
    END
  END O1[11]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 224.656 0.000 224.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 224.656 0.000 224.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 224.656 0.000 224.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 224.656 0.000 224.808 0.152 ;
    END
  END O1[10]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 224.352 0.000 224.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 224.352 0.000 224.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 224.352 0.000 224.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 224.352 0.000 224.504 0.152 ;
    END
  END O1[9]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 224.048 0.000 224.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 224.048 0.000 224.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 224.048 0.000 224.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 224.048 0.000 224.200 0.152 ;
    END
  END O1[8]

  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.832 0.000 222.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 222.832 0.000 222.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 222.832 0.000 222.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 222.832 0.000 222.984 0.152 ;
    END
  END I1[8]

  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.528 0.000 222.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 222.528 0.000 222.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 222.528 0.000 222.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 222.528 0.000 222.680 0.152 ;
    END
  END I1[9]

  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.224 0.000 222.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 222.224 0.000 222.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 222.224 0.000 222.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 222.224 0.000 222.376 0.152 ;
    END
  END I1[10]

  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 221.920 0.000 222.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 221.920 0.000 222.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 221.920 0.000 222.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 221.920 0.000 222.072 0.152 ;
    END
  END I1[11]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 220.704 0.000 220.856 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 220.704 0.000 220.856 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 220.704 0.000 220.856 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 220.704 0.000 220.856 0.152 ;
    END
  END O1[15]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 220.400 0.000 220.552 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 220.400 0.000 220.552 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 220.400 0.000 220.552 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 220.400 0.000 220.552 0.152 ;
    END
  END O1[14]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 220.096 0.000 220.248 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 220.096 0.000 220.248 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 220.096 0.000 220.248 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 220.096 0.000 220.248 0.152 ;
    END
  END O1[13]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.792 0.000 219.944 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 219.792 0.000 219.944 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 219.792 0.000 219.944 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 219.792 0.000 219.944 0.152 ;
    END
  END O1[12]

  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 218.576 0.000 218.728 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 218.576 0.000 218.728 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 218.576 0.000 218.728 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 218.576 0.000 218.728 0.152 ;
    END
  END I1[12]

  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 218.272 0.000 218.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 218.272 0.000 218.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 218.272 0.000 218.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 218.272 0.000 218.424 0.152 ;
    END
  END I1[13]

  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 217.968 0.000 218.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 217.968 0.000 218.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 217.968 0.000 218.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 217.968 0.000 218.120 0.152 ;
    END
  END I1[14]

  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 217.664 0.000 217.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 217.664 0.000 217.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 217.664 0.000 217.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 217.664 0.000 217.816 0.152 ;
    END
  END I1[15]

  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.448 0.000 216.600 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 216.448 0.000 216.600 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 216.448 0.000 216.600 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 216.448 0.000 216.600 0.152 ;
    END
  END O1[19]

  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.144 0.000 216.296 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 216.144 0.000 216.296 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 216.144 0.000 216.296 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 216.144 0.000 216.296 0.152 ;
    END
  END O1[18]

  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.840 0.000 215.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 215.840 0.000 215.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 215.840 0.000 215.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 215.840 0.000 215.992 0.152 ;
    END
  END O1[17]

  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.536 0.000 215.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 215.536 0.000 215.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 215.536 0.000 215.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 215.536 0.000 215.688 0.152 ;
    END
  END O1[16]

  PIN I1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 214.320 0.000 214.472 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 214.320 0.000 214.472 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 214.320 0.000 214.472 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 214.320 0.000 214.472 0.152 ;
    END
  END I1[16]

  PIN I1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 214.016 0.000 214.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 214.016 0.000 214.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 214.016 0.000 214.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 214.016 0.000 214.168 0.152 ;
    END
  END I1[17]

  PIN I1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 213.712 0.000 213.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 213.712 0.000 213.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 213.712 0.000 213.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 213.712 0.000 213.864 0.152 ;
    END
  END I1[18]

  PIN I1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 213.408 0.000 213.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 213.408 0.000 213.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 213.408 0.000 213.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 213.408 0.000 213.560 0.152 ;
    END
  END I1[19]

  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 212.192 0.000 212.344 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 212.192 0.000 212.344 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 212.192 0.000 212.344 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 212.192 0.000 212.344 0.152 ;
    END
  END O1[23]

  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.888 0.000 212.040 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 211.888 0.000 212.040 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 211.888 0.000 212.040 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 211.888 0.000 212.040 0.152 ;
    END
  END O1[22]

  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.584 0.000 211.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 211.584 0.000 211.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 211.584 0.000 211.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 211.584 0.000 211.736 0.152 ;
    END
  END O1[21]

  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.280 0.000 211.432 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 211.280 0.000 211.432 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 211.280 0.000 211.432 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 211.280 0.000 211.432 0.152 ;
    END
  END O1[20]

  PIN I1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 210.064 0.000 210.216 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 210.064 0.000 210.216 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 210.064 0.000 210.216 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 210.064 0.000 210.216 0.152 ;
    END
  END I1[20]

  PIN I1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 209.760 0.000 209.912 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 209.760 0.000 209.912 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 209.760 0.000 209.912 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 209.760 0.000 209.912 0.152 ;
    END
  END I1[21]

  PIN I1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 209.456 0.000 209.608 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 209.456 0.000 209.608 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 209.456 0.000 209.608 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 209.456 0.000 209.608 0.152 ;
    END
  END I1[22]

  PIN I1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 209.152 0.000 209.304 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 209.152 0.000 209.304 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 209.152 0.000 209.304 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 209.152 0.000 209.304 0.152 ;
    END
  END I1[23]

  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.936 0.000 208.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 207.936 0.000 208.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 207.936 0.000 208.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 207.936 0.000 208.088 0.152 ;
    END
  END O1[27]

  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.632 0.000 207.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 207.632 0.000 207.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 207.632 0.000 207.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 207.632 0.000 207.784 0.152 ;
    END
  END O1[26]

  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.328 0.000 207.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 207.328 0.000 207.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 207.328 0.000 207.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 207.328 0.000 207.480 0.152 ;
    END
  END O1[25]

  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.024 0.000 207.176 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 207.024 0.000 207.176 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 207.024 0.000 207.176 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 207.024 0.000 207.176 0.152 ;
    END
  END O1[24]

  PIN I1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.808 0.000 205.960 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.808 0.000 205.960 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.808 0.000 205.960 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.808 0.000 205.960 0.152 ;
    END
  END I1[24]

  PIN I1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.504 0.000 205.656 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.504 0.000 205.656 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.504 0.000 205.656 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.504 0.000 205.656 0.152 ;
    END
  END I1[25]

  PIN I1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.200 0.000 205.352 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.200 0.000 205.352 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.200 0.000 205.352 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.200 0.000 205.352 0.152 ;
    END
  END I1[26]

  PIN I1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.896 0.000 205.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 204.896 0.000 205.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 204.896 0.000 205.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 204.896 0.000 205.048 0.152 ;
    END
  END I1[27]

  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.680 0.000 203.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 203.680 0.000 203.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 203.680 0.000 203.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 203.680 0.000 203.832 0.152 ;
    END
  END O1[31]

  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.376 0.000 203.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 203.376 0.000 203.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 203.376 0.000 203.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 203.376 0.000 203.528 0.152 ;
    END
  END O1[30]

  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.072 0.000 203.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 203.072 0.000 203.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 203.072 0.000 203.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 203.072 0.000 203.224 0.152 ;
    END
  END O1[29]

  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 202.768 0.000 202.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 202.768 0.000 202.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 202.768 0.000 202.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 202.768 0.000 202.920 0.152 ;
    END
  END O1[28]

  PIN I1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 201.552 0.000 201.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 201.552 0.000 201.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 201.552 0.000 201.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 201.552 0.000 201.704 0.152 ;
    END
  END I1[28]

  PIN I1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 201.248 0.000 201.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 201.248 0.000 201.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 201.248 0.000 201.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 201.248 0.000 201.400 0.152 ;
    END
  END I1[29]

  PIN I1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 200.944 0.000 201.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 200.944 0.000 201.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 200.944 0.000 201.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 200.944 0.000 201.096 0.152 ;
    END
  END I1[30]

  PIN I1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 200.640 0.000 200.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 200.640 0.000 200.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 200.640 0.000 200.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 200.640 0.000 200.792 0.152 ;
    END
  END I1[31]

  PIN O1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 199.424 0.000 199.576 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 199.424 0.000 199.576 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 199.424 0.000 199.576 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 199.424 0.000 199.576 0.152 ;
    END
  END O1[35]

  PIN O1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 199.120 0.000 199.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 199.120 0.000 199.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 199.120 0.000 199.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 199.120 0.000 199.272 0.152 ;
    END
  END O1[34]

  PIN O1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 198.816 0.000 198.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 198.816 0.000 198.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 198.816 0.000 198.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 198.816 0.000 198.968 0.152 ;
    END
  END O1[33]

  PIN O1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 198.512 0.000 198.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 198.512 0.000 198.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 198.512 0.000 198.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 198.512 0.000 198.664 0.152 ;
    END
  END O1[32]

  PIN I1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 197.296 0.000 197.448 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.296 0.000 197.448 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.296 0.000 197.448 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 197.296 0.000 197.448 0.152 ;
    END
  END I1[32]

  PIN I1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.992 0.000 197.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 196.992 0.000 197.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 196.992 0.000 197.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 196.992 0.000 197.144 0.152 ;
    END
  END I1[33]

  PIN I1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.688 0.000 196.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 196.688 0.000 196.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 196.688 0.000 196.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 196.688 0.000 196.840 0.152 ;
    END
  END I1[34]

  PIN I1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.384 0.000 196.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 196.384 0.000 196.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 196.384 0.000 196.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 196.384 0.000 196.536 0.152 ;
    END
  END I1[35]

  PIN O1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 195.168 0.000 195.320 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 195.168 0.000 195.320 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 195.168 0.000 195.320 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 195.168 0.000 195.320 0.152 ;
    END
  END O1[39]

  PIN O1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.864 0.000 195.016 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 194.864 0.000 195.016 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 194.864 0.000 195.016 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 194.864 0.000 195.016 0.152 ;
    END
  END O1[38]

  PIN O1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.560 0.000 194.712 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 194.560 0.000 194.712 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 194.560 0.000 194.712 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 194.560 0.000 194.712 0.152 ;
    END
  END O1[37]

  PIN O1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.256 0.000 194.408 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 194.256 0.000 194.408 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 194.256 0.000 194.408 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 194.256 0.000 194.408 0.152 ;
    END
  END O1[36]

  PIN I1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 193.040 0.000 193.192 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 193.040 0.000 193.192 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 193.040 0.000 193.192 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 193.040 0.000 193.192 0.152 ;
    END
  END I1[36]

  PIN I1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.736 0.000 192.888 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 192.736 0.000 192.888 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 192.736 0.000 192.888 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 192.736 0.000 192.888 0.152 ;
    END
  END I1[37]

  PIN I1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.432 0.000 192.584 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 192.432 0.000 192.584 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 192.432 0.000 192.584 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 192.432 0.000 192.584 0.152 ;
    END
  END I1[38]

  PIN I1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.128 0.000 192.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 192.128 0.000 192.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 192.128 0.000 192.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 192.128 0.000 192.280 0.152 ;
    END
  END I1[39]

  PIN O1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.912 0.000 191.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 190.912 0.000 191.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 190.912 0.000 191.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.912 0.000 191.064 0.152 ;
    END
  END O1[43]

  PIN O1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
  END O1[42]

  PIN O1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.304 0.000 190.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 190.304 0.000 190.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 190.304 0.000 190.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.304 0.000 190.456 0.152 ;
    END
  END O1[41]

  PIN O1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.000 0.000 190.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 190.000 0.000 190.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 190.000 0.000 190.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.000 0.000 190.152 0.152 ;
    END
  END O1[40]

  PIN I1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 188.784 0.000 188.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 188.784 0.000 188.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 188.784 0.000 188.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 188.784 0.000 188.936 0.152 ;
    END
  END I1[40]

  PIN I1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 188.480 0.000 188.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 188.480 0.000 188.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 188.480 0.000 188.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 188.480 0.000 188.632 0.152 ;
    END
  END I1[41]

  PIN I1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 188.176 0.000 188.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 188.176 0.000 188.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 188.176 0.000 188.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 188.176 0.000 188.328 0.152 ;
    END
  END I1[42]

  PIN I1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 187.872 0.000 188.024 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 187.872 0.000 188.024 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 187.872 0.000 188.024 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 187.872 0.000 188.024 0.152 ;
    END
  END I1[43]

  PIN O1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.656 0.000 186.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 186.656 0.000 186.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 186.656 0.000 186.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 186.656 0.000 186.808 0.152 ;
    END
  END O1[47]

  PIN O1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.352 0.000 186.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 186.352 0.000 186.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 186.352 0.000 186.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 186.352 0.000 186.504 0.152 ;
    END
  END O1[46]

  PIN O1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.048 0.000 186.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 186.048 0.000 186.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 186.048 0.000 186.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 186.048 0.000 186.200 0.152 ;
    END
  END O1[45]

  PIN O1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 185.744 0.000 185.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 185.744 0.000 185.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 185.744 0.000 185.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 185.744 0.000 185.896 0.152 ;
    END
  END O1[44]

  PIN I1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 184.528 0.000 184.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 184.528 0.000 184.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 184.528 0.000 184.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 184.528 0.000 184.680 0.152 ;
    END
  END I1[44]

  PIN I1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 184.224 0.000 184.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 184.224 0.000 184.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 184.224 0.000 184.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 184.224 0.000 184.376 0.152 ;
    END
  END I1[45]

  PIN I1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.920 0.000 184.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 183.920 0.000 184.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 183.920 0.000 184.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 183.920 0.000 184.072 0.152 ;
    END
  END I1[46]

  PIN I1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.616 0.000 183.768 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 183.616 0.000 183.768 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 183.616 0.000 183.768 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 183.616 0.000 183.768 0.152 ;
    END
  END I1[47]

  PIN O1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 182.400 0.000 182.552 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 182.400 0.000 182.552 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 182.400 0.000 182.552 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 182.400 0.000 182.552 0.152 ;
    END
  END O1[51]

  PIN O1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 182.096 0.000 182.248 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 182.096 0.000 182.248 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 182.096 0.000 182.248 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 182.096 0.000 182.248 0.152 ;
    END
  END O1[50]

  PIN O1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 181.792 0.000 181.944 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 181.792 0.000 181.944 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 181.792 0.000 181.944 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 181.792 0.000 181.944 0.152 ;
    END
  END O1[49]

  PIN O1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 181.488 0.000 181.640 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 181.488 0.000 181.640 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 181.488 0.000 181.640 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 181.488 0.000 181.640 0.152 ;
    END
  END O1[48]

  PIN I1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 180.272 0.000 180.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 180.272 0.000 180.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 180.272 0.000 180.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 180.272 0.000 180.424 0.152 ;
    END
  END I1[48]

  PIN I1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.968 0.000 180.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 179.968 0.000 180.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 179.968 0.000 180.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 179.968 0.000 180.120 0.152 ;
    END
  END I1[49]

  PIN I1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.664 0.000 179.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 179.664 0.000 179.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 179.664 0.000 179.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 179.664 0.000 179.816 0.152 ;
    END
  END I1[50]

  PIN I1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.360 0.000 179.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 179.360 0.000 179.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 179.360 0.000 179.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 179.360 0.000 179.512 0.152 ;
    END
  END I1[51]

  PIN O1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.144 0.000 178.296 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 178.144 0.000 178.296 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 178.144 0.000 178.296 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 178.144 0.000 178.296 0.152 ;
    END
  END O1[55]

  PIN O1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.840 0.000 177.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 177.840 0.000 177.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 177.840 0.000 177.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 177.840 0.000 177.992 0.152 ;
    END
  END O1[54]

  PIN O1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.536 0.000 177.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 177.536 0.000 177.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 177.536 0.000 177.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 177.536 0.000 177.688 0.152 ;
    END
  END O1[53]

  PIN O1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.232 0.000 177.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 177.232 0.000 177.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 177.232 0.000 177.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 177.232 0.000 177.384 0.152 ;
    END
  END O1[52]

  PIN I1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.016 0.000 176.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 176.016 0.000 176.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 176.016 0.000 176.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 176.016 0.000 176.168 0.152 ;
    END
  END I1[52]

  PIN I1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.712 0.000 175.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 175.712 0.000 175.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 175.712 0.000 175.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.712 0.000 175.864 0.152 ;
    END
  END I1[53]

  PIN I1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.408 0.000 175.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 175.408 0.000 175.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 175.408 0.000 175.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.408 0.000 175.560 0.152 ;
    END
  END I1[54]

  PIN I1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.104 0.000 175.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 175.104 0.000 175.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 175.104 0.000 175.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.104 0.000 175.256 0.152 ;
    END
  END I1[55]

  PIN O1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 173.888 0.000 174.040 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 173.888 0.000 174.040 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 173.888 0.000 174.040 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 173.888 0.000 174.040 0.152 ;
    END
  END O1[59]

  PIN O1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 173.584 0.000 173.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 173.584 0.000 173.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 173.584 0.000 173.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 173.584 0.000 173.736 0.152 ;
    END
  END O1[58]

  PIN O1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 173.280 0.000 173.432 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 173.280 0.000 173.432 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 173.280 0.000 173.432 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 173.280 0.000 173.432 0.152 ;
    END
  END O1[57]

  PIN O1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 172.976 0.000 173.128 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 172.976 0.000 173.128 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 172.976 0.000 173.128 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 172.976 0.000 173.128 0.152 ;
    END
  END O1[56]

  PIN I1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.760 0.000 171.912 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 171.760 0.000 171.912 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 171.760 0.000 171.912 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 171.760 0.000 171.912 0.152 ;
    END
  END I1[56]

  PIN I1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.456 0.000 171.608 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 171.456 0.000 171.608 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 171.456 0.000 171.608 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 171.456 0.000 171.608 0.152 ;
    END
  END I1[57]

  PIN I1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.152 0.000 171.304 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 171.152 0.000 171.304 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 171.152 0.000 171.304 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 171.152 0.000 171.304 0.152 ;
    END
  END I1[58]

  PIN I1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.848 0.000 171.000 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 170.848 0.000 171.000 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 170.848 0.000 171.000 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 170.848 0.000 171.000 0.152 ;
    END
  END I1[59]

  PIN O1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 169.632 0.000 169.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 169.632 0.000 169.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 169.632 0.000 169.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 169.632 0.000 169.784 0.152 ;
    END
  END O1[63]

  PIN O1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 169.328 0.000 169.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 169.328 0.000 169.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 169.328 0.000 169.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 169.328 0.000 169.480 0.152 ;
    END
  END O1[62]

  PIN O1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 169.024 0.000 169.176 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 169.024 0.000 169.176 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 169.024 0.000 169.176 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 169.024 0.000 169.176 0.152 ;
    END
  END O1[61]

  PIN O1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.720 0.000 168.872 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 168.720 0.000 168.872 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 168.720 0.000 168.872 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 168.720 0.000 168.872 0.152 ;
    END
  END O1[60]

  PIN I1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.504 0.000 167.656 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 167.504 0.000 167.656 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 167.504 0.000 167.656 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 167.504 0.000 167.656 0.152 ;
    END
  END I1[60]

  PIN I1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.200 0.000 167.352 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 167.200 0.000 167.352 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 167.200 0.000 167.352 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 167.200 0.000 167.352 0.152 ;
    END
  END I1[61]

  PIN I1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.896 0.000 167.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 166.896 0.000 167.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 166.896 0.000 167.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 166.896 0.000 167.048 0.152 ;
    END
  END I1[62]

  PIN I1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 166.592 0.000 166.744 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 166.592 0.000 166.744 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 166.592 0.000 166.744 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 166.592 0.000 166.744 0.152 ;
    END
  END I1[63]

  PIN O1[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.376 0.000 165.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 165.376 0.000 165.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 165.376 0.000 165.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 165.376 0.000 165.528 0.152 ;
    END
  END O1[67]

  PIN O1[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.072 0.000 165.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 165.072 0.000 165.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 165.072 0.000 165.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 165.072 0.000 165.224 0.152 ;
    END
  END O1[66]

  PIN O1[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.768 0.000 164.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 164.768 0.000 164.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 164.768 0.000 164.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 164.768 0.000 164.920 0.152 ;
    END
  END O1[65]

  PIN O1[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.464 0.000 164.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 164.464 0.000 164.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 164.464 0.000 164.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 164.464 0.000 164.616 0.152 ;
    END
  END O1[64]

  PIN I1[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 163.248 0.000 163.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 163.248 0.000 163.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 163.248 0.000 163.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 163.248 0.000 163.400 0.152 ;
    END
  END I1[64]

  PIN I1[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.944 0.000 163.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 162.944 0.000 163.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 162.944 0.000 163.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 162.944 0.000 163.096 0.152 ;
    END
  END I1[65]

  PIN I1[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.640 0.000 162.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 162.640 0.000 162.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 162.640 0.000 162.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 162.640 0.000 162.792 0.152 ;
    END
  END I1[66]

  PIN I1[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.336 0.000 162.488 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 162.336 0.000 162.488 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 162.336 0.000 162.488 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 162.336 0.000 162.488 0.152 ;
    END
  END I1[67]

  PIN O1[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.120 0.000 161.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 161.120 0.000 161.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 161.120 0.000 161.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.120 0.000 161.272 0.152 ;
    END
  END O1[71]

  PIN O1[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.816 0.000 160.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 160.816 0.000 160.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 160.816 0.000 160.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 160.816 0.000 160.968 0.152 ;
    END
  END O1[70]

  PIN O1[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.512 0.000 160.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 160.512 0.000 160.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 160.512 0.000 160.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 160.512 0.000 160.664 0.152 ;
    END
  END O1[69]

  PIN O1[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.208 0.000 160.360 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 160.208 0.000 160.360 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 160.208 0.000 160.360 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 160.208 0.000 160.360 0.152 ;
    END
  END O1[68]

  PIN I1[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.992 0.000 159.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 158.992 0.000 159.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 158.992 0.000 159.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 158.992 0.000 159.144 0.152 ;
    END
  END I1[68]

  PIN I1[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.688 0.000 158.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 158.688 0.000 158.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 158.688 0.000 158.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 158.688 0.000 158.840 0.152 ;
    END
  END I1[69]

  PIN I1[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.384 0.000 158.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 158.384 0.000 158.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 158.384 0.000 158.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 158.384 0.000 158.536 0.152 ;
    END
  END I1[70]

  PIN I1[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.080 0.000 158.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 158.080 0.000 158.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 158.080 0.000 158.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 158.080 0.000 158.232 0.152 ;
    END
  END I1[71]

  PIN O1[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.864 0.000 157.016 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 156.864 0.000 157.016 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 156.864 0.000 157.016 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 156.864 0.000 157.016 0.152 ;
    END
  END O1[75]

  PIN O1[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.560 0.000 156.712 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 156.560 0.000 156.712 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 156.560 0.000 156.712 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 156.560 0.000 156.712 0.152 ;
    END
  END O1[74]

  PIN O1[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.256 0.000 156.408 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 156.256 0.000 156.408 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 156.256 0.000 156.408 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 156.256 0.000 156.408 0.152 ;
    END
  END O1[73]

  PIN O1[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.952 0.000 156.104 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 155.952 0.000 156.104 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 155.952 0.000 156.104 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 155.952 0.000 156.104 0.152 ;
    END
  END O1[72]

  PIN I1[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.736 0.000 154.888 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.736 0.000 154.888 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.736 0.000 154.888 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 154.736 0.000 154.888 0.152 ;
    END
  END I1[72]

  PIN I1[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.432 0.000 154.584 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.432 0.000 154.584 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.432 0.000 154.584 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 154.432 0.000 154.584 0.152 ;
    END
  END I1[73]

  PIN I1[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
  END I1[74]

  PIN I1[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
  END I1[75]

  PIN O1[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.608 0.000 152.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 152.608 0.000 152.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 152.608 0.000 152.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 152.608 0.000 152.760 0.152 ;
    END
  END O1[79]

  PIN O1[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.304 0.000 152.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 152.304 0.000 152.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 152.304 0.000 152.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 152.304 0.000 152.456 0.152 ;
    END
  END O1[78]

  PIN O1[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.000 0.000 152.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 152.000 0.000 152.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 152.000 0.000 152.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 152.000 0.000 152.152 0.152 ;
    END
  END O1[77]

  PIN O1[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 151.696 0.000 151.848 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 151.696 0.000 151.848 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 151.696 0.000 151.848 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 151.696 0.000 151.848 0.152 ;
    END
  END O1[76]

  PIN I1[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.480 0.000 150.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.480 0.000 150.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.480 0.000 150.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 150.480 0.000 150.632 0.152 ;
    END
  END I1[76]

  PIN I1[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.176 0.000 150.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.176 0.000 150.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.176 0.000 150.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 150.176 0.000 150.328 0.152 ;
    END
  END I1[77]

  PIN I1[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.872 0.000 150.024 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 149.872 0.000 150.024 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 149.872 0.000 150.024 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 149.872 0.000 150.024 0.152 ;
    END
  END I1[78]

  PIN I1[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.568 0.000 149.720 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 149.568 0.000 149.720 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 149.568 0.000 149.720 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 149.568 0.000 149.720 0.152 ;
    END
  END I1[79]

  PIN O1[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.352 0.000 148.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.352 0.000 148.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.352 0.000 148.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.352 0.000 148.504 0.152 ;
    END
  END O1[83]

  PIN O1[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.048 0.000 148.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.048 0.000 148.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.048 0.000 148.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.048 0.000 148.200 0.152 ;
    END
  END O1[82]

  PIN O1[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.744 0.000 147.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 147.744 0.000 147.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 147.744 0.000 147.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 147.744 0.000 147.896 0.152 ;
    END
  END O1[81]

  PIN O1[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.440 0.000 147.592 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 147.440 0.000 147.592 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 147.440 0.000 147.592 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 147.440 0.000 147.592 0.152 ;
    END
  END O1[80]

  PIN I1[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.224 0.000 146.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 146.224 0.000 146.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 146.224 0.000 146.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.224 0.000 146.376 0.152 ;
    END
  END I1[80]

  PIN I1[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.920 0.000 146.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 145.920 0.000 146.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 145.920 0.000 146.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.920 0.000 146.072 0.152 ;
    END
  END I1[81]

  PIN I1[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.616 0.000 145.768 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 145.616 0.000 145.768 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 145.616 0.000 145.768 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.616 0.000 145.768 0.152 ;
    END
  END I1[82]

  PIN I1[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.312 0.000 145.464 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 145.312 0.000 145.464 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 145.312 0.000 145.464 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.312 0.000 145.464 0.152 ;
    END
  END I1[83]

  PIN O1[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.096 0.000 144.248 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 144.096 0.000 144.248 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 144.096 0.000 144.248 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 144.096 0.000 144.248 0.152 ;
    END
  END O1[87]

  PIN O1[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.792 0.000 143.944 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 143.792 0.000 143.944 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 143.792 0.000 143.944 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 143.792 0.000 143.944 0.152 ;
    END
  END O1[86]

  PIN O1[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.488 0.000 143.640 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 143.488 0.000 143.640 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 143.488 0.000 143.640 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 143.488 0.000 143.640 0.152 ;
    END
  END O1[85]

  PIN O1[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.184 0.000 143.336 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 143.184 0.000 143.336 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 143.184 0.000 143.336 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 143.184 0.000 143.336 0.152 ;
    END
  END O1[84]

  PIN I1[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.968 0.000 142.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 141.968 0.000 142.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.968 0.000 142.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.968 0.000 142.120 0.152 ;
    END
  END I1[84]

  PIN I1[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.664 0.000 141.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 141.664 0.000 141.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.664 0.000 141.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.664 0.000 141.816 0.152 ;
    END
  END I1[85]

  PIN I1[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.360 0.000 141.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 141.360 0.000 141.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.360 0.000 141.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.360 0.000 141.512 0.152 ;
    END
  END I1[86]

  PIN I1[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.056 0.000 141.208 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 141.056 0.000 141.208 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.056 0.000 141.208 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.056 0.000 141.208 0.152 ;
    END
  END I1[87]

  PIN O1[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.840 0.000 139.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 139.840 0.000 139.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 139.840 0.000 139.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 139.840 0.000 139.992 0.152 ;
    END
  END O1[91]

  PIN O1[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.536 0.000 139.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 139.536 0.000 139.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 139.536 0.000 139.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 139.536 0.000 139.688 0.152 ;
    END
  END O1[90]

  PIN O1[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.232 0.000 139.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 139.232 0.000 139.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 139.232 0.000 139.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 139.232 0.000 139.384 0.152 ;
    END
  END O1[89]

  PIN O1[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.928 0.000 139.080 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 138.928 0.000 139.080 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 138.928 0.000 139.080 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 138.928 0.000 139.080 0.152 ;
    END
  END O1[88]

  PIN I1[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.712 0.000 137.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 137.712 0.000 137.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 137.712 0.000 137.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 137.712 0.000 137.864 0.152 ;
    END
  END I1[88]

  PIN I1[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.408 0.000 137.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 137.408 0.000 137.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 137.408 0.000 137.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 137.408 0.000 137.560 0.152 ;
    END
  END I1[89]

  PIN I1[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.104 0.000 137.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 137.104 0.000 137.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 137.104 0.000 137.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 137.104 0.000 137.256 0.152 ;
    END
  END I1[90]

  PIN I1[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.800 0.000 136.952 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 136.800 0.000 136.952 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 136.800 0.000 136.952 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 136.800 0.000 136.952 0.152 ;
    END
  END I1[91]

  PIN O1[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.584 0.000 135.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 135.584 0.000 135.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 135.584 0.000 135.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 135.584 0.000 135.736 0.152 ;
    END
  END O1[95]

  PIN O1[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.280 0.000 135.432 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 135.280 0.000 135.432 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 135.280 0.000 135.432 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 135.280 0.000 135.432 0.152 ;
    END
  END O1[94]

  PIN O1[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.976 0.000 135.128 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 134.976 0.000 135.128 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 134.976 0.000 135.128 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.976 0.000 135.128 0.152 ;
    END
  END O1[93]

  PIN O1[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.672 0.000 134.824 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 134.672 0.000 134.824 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 134.672 0.000 134.824 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.672 0.000 134.824 0.152 ;
    END
  END O1[92]

  PIN I1[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.456 0.000 133.608 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 133.456 0.000 133.608 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 133.456 0.000 133.608 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 133.456 0.000 133.608 0.152 ;
    END
  END I1[92]

  PIN I1[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.152 0.000 133.304 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 133.152 0.000 133.304 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 133.152 0.000 133.304 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 133.152 0.000 133.304 0.152 ;
    END
  END I1[93]

  PIN I1[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.848 0.000 133.000 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.848 0.000 133.000 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.848 0.000 133.000 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 132.848 0.000 133.000 0.152 ;
    END
  END I1[94]

  PIN I1[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.544 0.000 132.696 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.544 0.000 132.696 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.544 0.000 132.696 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 132.544 0.000 132.696 0.152 ;
    END
  END I1[95]

  PIN O1[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.328 0.000 131.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.328 0.000 131.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.328 0.000 131.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.328 0.000 131.480 0.152 ;
    END
  END O1[99]

  PIN O1[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.024 0.000 131.176 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.024 0.000 131.176 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.024 0.000 131.176 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.024 0.000 131.176 0.152 ;
    END
  END O1[98]

  PIN O1[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.720 0.000 130.872 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 130.720 0.000 130.872 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 130.720 0.000 130.872 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.720 0.000 130.872 0.152 ;
    END
  END O1[97]

  PIN O1[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.416 0.000 130.568 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 130.416 0.000 130.568 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 130.416 0.000 130.568 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.416 0.000 130.568 0.152 ;
    END
  END O1[96]

  PIN I1[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.200 0.000 129.352 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 129.200 0.000 129.352 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 129.200 0.000 129.352 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.200 0.000 129.352 0.152 ;
    END
  END I1[96]

  PIN I1[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.896 0.000 129.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 128.896 0.000 129.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 128.896 0.000 129.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.896 0.000 129.048 0.152 ;
    END
  END I1[97]

  PIN I1[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.592 0.000 128.744 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 128.592 0.000 128.744 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 128.592 0.000 128.744 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.592 0.000 128.744 0.152 ;
    END
  END I1[98]

  PIN I1[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.288 0.000 128.440 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 128.288 0.000 128.440 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 128.288 0.000 128.440 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.288 0.000 128.440 0.152 ;
    END
  END I1[99]

  PIN O1[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.072 0.000 127.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 127.072 0.000 127.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 127.072 0.000 127.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.072 0.000 127.224 0.152 ;
    END
  END O1[103]

  PIN O1[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.768 0.000 126.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 126.768 0.000 126.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 126.768 0.000 126.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.768 0.000 126.920 0.152 ;
    END
  END O1[102]

  PIN O1[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.464 0.000 126.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 126.464 0.000 126.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 126.464 0.000 126.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.464 0.000 126.616 0.152 ;
    END
  END O1[101]

  PIN O1[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.160 0.000 126.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 126.160 0.000 126.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 126.160 0.000 126.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.160 0.000 126.312 0.152 ;
    END
  END O1[100]

  PIN I1[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.944 0.000 125.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 124.944 0.000 125.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 124.944 0.000 125.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.944 0.000 125.096 0.152 ;
    END
  END I1[100]

  PIN I1[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.640 0.000 124.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 124.640 0.000 124.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 124.640 0.000 124.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.640 0.000 124.792 0.152 ;
    END
  END I1[101]

  PIN I1[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.336 0.000 124.488 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 124.336 0.000 124.488 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 124.336 0.000 124.488 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.336 0.000 124.488 0.152 ;
    END
  END I1[102]

  PIN I1[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.032 0.000 124.184 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 124.032 0.000 124.184 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 124.032 0.000 124.184 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.032 0.000 124.184 0.152 ;
    END
  END I1[103]

  PIN O1[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.816 0.000 122.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 122.816 0.000 122.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 122.816 0.000 122.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.816 0.000 122.968 0.152 ;
    END
  END O1[107]

  PIN O1[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.512 0.000 122.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 122.512 0.000 122.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 122.512 0.000 122.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.512 0.000 122.664 0.152 ;
    END
  END O1[106]

  PIN O1[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.208 0.000 122.360 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 122.208 0.000 122.360 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 122.208 0.000 122.360 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.208 0.000 122.360 0.152 ;
    END
  END O1[105]

  PIN O1[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.904 0.000 122.056 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 121.904 0.000 122.056 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 121.904 0.000 122.056 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.904 0.000 122.056 0.152 ;
    END
  END O1[104]

  PIN I1[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.688 0.000 120.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.688 0.000 120.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.688 0.000 120.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.688 0.000 120.840 0.152 ;
    END
  END I1[104]

  PIN I1[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.384 0.000 120.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.384 0.000 120.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.384 0.000 120.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.384 0.000 120.536 0.152 ;
    END
  END I1[105]

  PIN I1[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.080 0.000 120.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.080 0.000 120.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.080 0.000 120.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.080 0.000 120.232 0.152 ;
    END
  END I1[106]

  PIN I1[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.776 0.000 119.928 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 119.776 0.000 119.928 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 119.776 0.000 119.928 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.776 0.000 119.928 0.152 ;
    END
  END I1[107]

  PIN O1[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.560 0.000 118.712 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 118.560 0.000 118.712 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 118.560 0.000 118.712 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.560 0.000 118.712 0.152 ;
    END
  END O1[111]

  PIN O1[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.256 0.000 118.408 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 118.256 0.000 118.408 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 118.256 0.000 118.408 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.256 0.000 118.408 0.152 ;
    END
  END O1[110]

  PIN O1[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.952 0.000 118.104 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 117.952 0.000 118.104 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 117.952 0.000 118.104 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.952 0.000 118.104 0.152 ;
    END
  END O1[109]

  PIN O1[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.648 0.000 117.800 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 117.648 0.000 117.800 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 117.648 0.000 117.800 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.648 0.000 117.800 0.152 ;
    END
  END O1[108]

  PIN I1[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.432 0.000 116.584 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 116.432 0.000 116.584 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 116.432 0.000 116.584 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.432 0.000 116.584 0.152 ;
    END
  END I1[108]

  PIN I1[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.128 0.000 116.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 116.128 0.000 116.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 116.128 0.000 116.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.128 0.000 116.280 0.152 ;
    END
  END I1[109]

  PIN I1[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.824 0.000 115.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 115.824 0.000 115.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 115.824 0.000 115.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.824 0.000 115.976 0.152 ;
    END
  END I1[110]

  PIN I1[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.520 0.000 115.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 115.520 0.000 115.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 115.520 0.000 115.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.520 0.000 115.672 0.152 ;
    END
  END I1[111]

  PIN O1[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.304 0.000 114.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 114.304 0.000 114.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 114.304 0.000 114.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.304 0.000 114.456 0.152 ;
    END
  END O1[115]

  PIN O1[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.000 0.000 114.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 114.000 0.000 114.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 114.000 0.000 114.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.000 0.000 114.152 0.152 ;
    END
  END O1[114]

  PIN O1[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.696 0.000 113.848 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 113.696 0.000 113.848 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 113.696 0.000 113.848 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.696 0.000 113.848 0.152 ;
    END
  END O1[113]

  PIN O1[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.392 0.000 113.544 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 113.392 0.000 113.544 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 113.392 0.000 113.544 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.392 0.000 113.544 0.152 ;
    END
  END O1[112]

  PIN I1[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.176 0.000 112.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 112.176 0.000 112.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.176 0.000 112.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.176 0.000 112.328 0.152 ;
    END
  END I1[112]

  PIN I1[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.872 0.000 112.024 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 111.872 0.000 112.024 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 111.872 0.000 112.024 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.872 0.000 112.024 0.152 ;
    END
  END I1[113]

  PIN I1[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.568 0.000 111.720 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 111.568 0.000 111.720 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 111.568 0.000 111.720 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.568 0.000 111.720 0.152 ;
    END
  END I1[114]

  PIN I1[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.264 0.000 111.416 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 111.264 0.000 111.416 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 111.264 0.000 111.416 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.264 0.000 111.416 0.152 ;
    END
  END I1[115]

  PIN O1[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
  END O1[119]

  PIN O1[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.744 0.000 109.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.744 0.000 109.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.744 0.000 109.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.744 0.000 109.896 0.152 ;
    END
  END O1[118]

  PIN O1[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.440 0.000 109.592 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.440 0.000 109.592 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.440 0.000 109.592 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.440 0.000 109.592 0.152 ;
    END
  END O1[117]

  PIN O1[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.136 0.000 109.288 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.136 0.000 109.288 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.136 0.000 109.288 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.136 0.000 109.288 0.152 ;
    END
  END O1[116]

  PIN I1[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.920 0.000 108.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.920 0.000 108.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.920 0.000 108.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.920 0.000 108.072 0.152 ;
    END
  END I1[116]

  PIN I1[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.616 0.000 107.768 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.616 0.000 107.768 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.616 0.000 107.768 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.616 0.000 107.768 0.152 ;
    END
  END I1[117]

  PIN I1[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.312 0.000 107.464 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.312 0.000 107.464 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.312 0.000 107.464 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.312 0.000 107.464 0.152 ;
    END
  END I1[118]

  PIN I1[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.008 0.000 107.160 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.008 0.000 107.160 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.008 0.000 107.160 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.008 0.000 107.160 0.152 ;
    END
  END I1[119]

  PIN O1[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.792 0.000 105.944 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.792 0.000 105.944 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.792 0.000 105.944 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.792 0.000 105.944 0.152 ;
    END
  END O1[123]

  PIN O1[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.488 0.000 105.640 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.488 0.000 105.640 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.488 0.000 105.640 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.488 0.000 105.640 0.152 ;
    END
  END O1[122]

  PIN O1[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.184 0.000 105.336 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.184 0.000 105.336 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.184 0.000 105.336 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.184 0.000 105.336 0.152 ;
    END
  END O1[121]

  PIN O1[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.880 0.000 105.032 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.880 0.000 105.032 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.880 0.000 105.032 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.880 0.000 105.032 0.152 ;
    END
  END O1[120]

  PIN I1[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.664 0.000 103.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.664 0.000 103.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.664 0.000 103.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.664 0.000 103.816 0.152 ;
    END
  END I1[120]

  PIN I1[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.360 0.000 103.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.360 0.000 103.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.360 0.000 103.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.360 0.000 103.512 0.152 ;
    END
  END I1[121]

  PIN I1[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.056 0.000 103.208 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.056 0.000 103.208 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.056 0.000 103.208 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.056 0.000 103.208 0.152 ;
    END
  END I1[122]

  PIN I1[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.752 0.000 102.904 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.752 0.000 102.904 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.752 0.000 102.904 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.752 0.000 102.904 0.152 ;
    END
  END I1[123]

  PIN O1[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.536 0.000 101.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.536 0.000 101.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.536 0.000 101.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.536 0.000 101.688 0.152 ;
    END
  END O1[127]

  PIN O1[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.232 0.000 101.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.232 0.000 101.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.232 0.000 101.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.232 0.000 101.384 0.152 ;
    END
  END O1[126]

  PIN O1[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.928 0.000 101.080 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.928 0.000 101.080 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.928 0.000 101.080 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.928 0.000 101.080 0.152 ;
    END
  END O1[125]

  PIN O1[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.624 0.000 100.776 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.624 0.000 100.776 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.624 0.000 100.776 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.624 0.000 100.776 0.152 ;
    END
  END O1[124]

  PIN I1[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.408 0.000 99.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.408 0.000 99.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.408 0.000 99.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.408 0.000 99.560 0.152 ;
    END
  END I1[124]

  PIN I1[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.104 0.000 99.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.104 0.000 99.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.104 0.000 99.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.104 0.000 99.256 0.152 ;
    END
  END I1[125]

  PIN I1[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.800 0.000 98.952 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.800 0.000 98.952 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.800 0.000 98.952 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.800 0.000 98.952 0.152 ;
    END
  END I1[126]

  PIN I1[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.496 0.000 98.648 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.496 0.000 98.648 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.496 0.000 98.648 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.496 0.000 98.648 0.152 ;
    END
  END I1[127]

  PIN O1[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.280 0.000 97.432 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.280 0.000 97.432 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.280 0.000 97.432 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.280 0.000 97.432 0.152 ;
    END
  END O1[131]

  PIN O1[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.976 0.000 97.128 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.976 0.000 97.128 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.976 0.000 97.128 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.976 0.000 97.128 0.152 ;
    END
  END O1[130]

  PIN O1[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.672 0.000 96.824 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.672 0.000 96.824 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.672 0.000 96.824 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.672 0.000 96.824 0.152 ;
    END
  END O1[129]

  PIN O1[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.368 0.000 96.520 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.368 0.000 96.520 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.368 0.000 96.520 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.368 0.000 96.520 0.152 ;
    END
  END O1[128]

  PIN I1[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.152 0.000 95.304 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.152 0.000 95.304 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.152 0.000 95.304 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.152 0.000 95.304 0.152 ;
    END
  END I1[128]

  PIN I1[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.848 0.000 95.000 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.848 0.000 95.000 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.848 0.000 95.000 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.848 0.000 95.000 0.152 ;
    END
  END I1[129]

  PIN I1[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.544 0.000 94.696 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.544 0.000 94.696 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.544 0.000 94.696 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.544 0.000 94.696 0.152 ;
    END
  END I1[130]

  PIN I1[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.240 0.000 94.392 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.240 0.000 94.392 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.240 0.000 94.392 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.240 0.000 94.392 0.152 ;
    END
  END I1[131]

  PIN O1[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
  END O1[135]

  PIN O1[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.720 0.000 92.872 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.720 0.000 92.872 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.720 0.000 92.872 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.720 0.000 92.872 0.152 ;
    END
  END O1[134]

  PIN O1[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.416 0.000 92.568 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.416 0.000 92.568 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.416 0.000 92.568 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.416 0.000 92.568 0.152 ;
    END
  END O1[133]

  PIN O1[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.112 0.000 92.264 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.112 0.000 92.264 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.112 0.000 92.264 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.112 0.000 92.264 0.152 ;
    END
  END O1[132]

  PIN I1[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.896 0.000 91.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.896 0.000 91.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.896 0.000 91.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.896 0.000 91.048 0.152 ;
    END
  END I1[132]

  PIN I1[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.592 0.000 90.744 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.592 0.000 90.744 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.592 0.000 90.744 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.592 0.000 90.744 0.152 ;
    END
  END I1[133]

  PIN I1[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.288 0.000 90.440 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.288 0.000 90.440 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.288 0.000 90.440 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.288 0.000 90.440 0.152 ;
    END
  END I1[134]

  PIN I1[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.984 0.000 90.136 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.984 0.000 90.136 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.984 0.000 90.136 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.984 0.000 90.136 0.152 ;
    END
  END I1[135]

  PIN O1[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
  END O1[139]

  PIN O1[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
  END O1[138]

  PIN O1[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
  END O1[137]

  PIN O1[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
  END O1[136]

  PIN I1[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.640 0.000 86.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.640 0.000 86.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.640 0.000 86.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.640 0.000 86.792 0.152 ;
    END
  END I1[136]

  PIN I1[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.336 0.000 86.488 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.336 0.000 86.488 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.336 0.000 86.488 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.336 0.000 86.488 0.152 ;
    END
  END I1[137]

  PIN I1[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.032 0.000 86.184 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.032 0.000 86.184 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.032 0.000 86.184 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.032 0.000 86.184 0.152 ;
    END
  END I1[138]

  PIN I1[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.728 0.000 85.880 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.728 0.000 85.880 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.728 0.000 85.880 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.728 0.000 85.880 0.152 ;
    END
  END I1[139]

  PIN O1[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.512 0.000 84.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.512 0.000 84.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.512 0.000 84.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.512 0.000 84.664 0.152 ;
    END
  END O1[143]

  PIN O1[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.208 0.000 84.360 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.208 0.000 84.360 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.208 0.000 84.360 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.208 0.000 84.360 0.152 ;
    END
  END O1[142]

  PIN O1[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.904 0.000 84.056 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.904 0.000 84.056 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.904 0.000 84.056 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.904 0.000 84.056 0.152 ;
    END
  END O1[141]

  PIN O1[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.600 0.000 83.752 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.600 0.000 83.752 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.600 0.000 83.752 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.600 0.000 83.752 0.152 ;
    END
  END O1[140]

  PIN I1[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
  END I1[140]

  PIN I1[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.080 0.000 82.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.080 0.000 82.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.080 0.000 82.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.080 0.000 82.232 0.152 ;
    END
  END I1[141]

  PIN I1[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.776 0.000 81.928 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.776 0.000 81.928 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.776 0.000 81.928 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.776 0.000 81.928 0.152 ;
    END
  END I1[142]

  PIN I1[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.472 0.000 81.624 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.472 0.000 81.624 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.472 0.000 81.624 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.472 0.000 81.624 0.152 ;
    END
  END I1[143]

  PIN O1[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.256 0.000 80.408 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.256 0.000 80.408 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.256 0.000 80.408 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.256 0.000 80.408 0.152 ;
    END
  END O1[147]

  PIN O1[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.952 0.000 80.104 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.952 0.000 80.104 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.952 0.000 80.104 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.952 0.000 80.104 0.152 ;
    END
  END O1[146]

  PIN O1[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.648 0.000 79.800 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.648 0.000 79.800 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.648 0.000 79.800 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.648 0.000 79.800 0.152 ;
    END
  END O1[145]

  PIN O1[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.344 0.000 79.496 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.344 0.000 79.496 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.344 0.000 79.496 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.344 0.000 79.496 0.152 ;
    END
  END O1[144]

  PIN I1[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.128 0.000 78.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.128 0.000 78.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.128 0.000 78.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.128 0.000 78.280 0.152 ;
    END
  END I1[144]

  PIN I1[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.824 0.000 77.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.824 0.000 77.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.824 0.000 77.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.824 0.000 77.976 0.152 ;
    END
  END I1[145]

  PIN I1[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.520 0.000 77.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.520 0.000 77.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.520 0.000 77.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.520 0.000 77.672 0.152 ;
    END
  END I1[146]

  PIN I1[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.216 0.000 77.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.216 0.000 77.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.216 0.000 77.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.216 0.000 77.368 0.152 ;
    END
  END I1[147]

  PIN O1[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.000 0.000 76.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.000 0.000 76.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.000 0.000 76.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.000 0.000 76.152 0.152 ;
    END
  END O1[151]

  PIN O1[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.696 0.000 75.848 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.696 0.000 75.848 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.696 0.000 75.848 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.696 0.000 75.848 0.152 ;
    END
  END O1[150]

  PIN O1[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.392 0.000 75.544 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.392 0.000 75.544 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.392 0.000 75.544 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.392 0.000 75.544 0.152 ;
    END
  END O1[149]

  PIN O1[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.088 0.000 75.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.088 0.000 75.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.088 0.000 75.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.088 0.000 75.240 0.152 ;
    END
  END O1[148]

  PIN I1[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.872 0.000 74.024 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.872 0.000 74.024 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.872 0.000 74.024 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.872 0.000 74.024 0.152 ;
    END
  END I1[148]

  PIN I1[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.568 0.000 73.720 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.568 0.000 73.720 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.568 0.000 73.720 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.568 0.000 73.720 0.152 ;
    END
  END I1[149]

  PIN I1[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.264 0.000 73.416 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.264 0.000 73.416 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.264 0.000 73.416 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.264 0.000 73.416 0.152 ;
    END
  END I1[150]

  PIN I1[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.960 0.000 73.112 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.960 0.000 73.112 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.960 0.000 73.112 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.960 0.000 73.112 0.152 ;
    END
  END I1[151]

  PIN O1[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
  END O1[155]

  PIN O1[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.440 0.000 71.592 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.440 0.000 71.592 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.440 0.000 71.592 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.440 0.000 71.592 0.152 ;
    END
  END O1[154]

  PIN O1[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.136 0.000 71.288 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.136 0.000 71.288 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.136 0.000 71.288 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.136 0.000 71.288 0.152 ;
    END
  END O1[153]

  PIN O1[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.832 0.000 70.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.832 0.000 70.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.832 0.000 70.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.832 0.000 70.984 0.152 ;
    END
  END O1[152]

  PIN I1[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.616 0.000 69.768 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.616 0.000 69.768 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.616 0.000 69.768 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.616 0.000 69.768 0.152 ;
    END
  END I1[152]

  PIN I1[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.312 0.000 69.464 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.312 0.000 69.464 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.312 0.000 69.464 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.312 0.000 69.464 0.152 ;
    END
  END I1[153]

  PIN I1[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.008 0.000 69.160 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.008 0.000 69.160 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.008 0.000 69.160 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.008 0.000 69.160 0.152 ;
    END
  END I1[154]

  PIN I1[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.704 0.000 68.856 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.704 0.000 68.856 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.704 0.000 68.856 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.704 0.000 68.856 0.152 ;
    END
  END I1[155]

  PIN O1[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.488 0.000 67.640 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.488 0.000 67.640 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.488 0.000 67.640 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.488 0.000 67.640 0.152 ;
    END
  END O1[159]

  PIN O1[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.184 0.000 67.336 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.184 0.000 67.336 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.184 0.000 67.336 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.184 0.000 67.336 0.152 ;
    END
  END O1[158]

  PIN O1[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.880 0.000 67.032 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.880 0.000 67.032 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.880 0.000 67.032 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.880 0.000 67.032 0.152 ;
    END
  END O1[157]

  PIN O1[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.576 0.000 66.728 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.576 0.000 66.728 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.576 0.000 66.728 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.576 0.000 66.728 0.152 ;
    END
  END O1[156]

  PIN I1[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.360 0.000 65.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.360 0.000 65.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.360 0.000 65.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.360 0.000 65.512 0.152 ;
    END
  END I1[156]

  PIN I1[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.056 0.000 65.208 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.056 0.000 65.208 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.056 0.000 65.208 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.056 0.000 65.208 0.152 ;
    END
  END I1[157]

  PIN I1[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.752 0.000 64.904 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.752 0.000 64.904 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.752 0.000 64.904 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.752 0.000 64.904 0.152 ;
    END
  END I1[158]

  PIN I1[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.448 0.000 64.600 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.448 0.000 64.600 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.448 0.000 64.600 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.448 0.000 64.600 0.152 ;
    END
  END I1[159]

  PIN O1[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.232 0.000 63.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.232 0.000 63.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.232 0.000 63.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.232 0.000 63.384 0.152 ;
    END
  END O1[163]

  PIN O1[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.928 0.000 63.080 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.928 0.000 63.080 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.928 0.000 63.080 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.928 0.000 63.080 0.152 ;
    END
  END O1[162]

  PIN O1[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.624 0.000 62.776 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.624 0.000 62.776 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.624 0.000 62.776 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.624 0.000 62.776 0.152 ;
    END
  END O1[161]

  PIN O1[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.320 0.000 62.472 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.320 0.000 62.472 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.320 0.000 62.472 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.320 0.000 62.472 0.152 ;
    END
  END O1[160]

  PIN I1[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.104 0.000 61.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.104 0.000 61.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.104 0.000 61.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.104 0.000 61.256 0.152 ;
    END
  END I1[160]

  PIN I1[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.800 0.000 60.952 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.800 0.000 60.952 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.800 0.000 60.952 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.800 0.000 60.952 0.152 ;
    END
  END I1[161]

  PIN I1[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.496 0.000 60.648 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.496 0.000 60.648 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.496 0.000 60.648 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.496 0.000 60.648 0.152 ;
    END
  END I1[162]

  PIN I1[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.192 0.000 60.344 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.192 0.000 60.344 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.192 0.000 60.344 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.192 0.000 60.344 0.152 ;
    END
  END I1[163]

  PIN O1[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.976 0.000 59.128 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.976 0.000 59.128 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.976 0.000 59.128 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.976 0.000 59.128 0.152 ;
    END
  END O1[167]

  PIN O1[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.672 0.000 58.824 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.672 0.000 58.824 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.672 0.000 58.824 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.672 0.000 58.824 0.152 ;
    END
  END O1[166]

  PIN O1[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.368 0.000 58.520 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.368 0.000 58.520 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.368 0.000 58.520 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.368 0.000 58.520 0.152 ;
    END
  END O1[165]

  PIN O1[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.064 0.000 58.216 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.064 0.000 58.216 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.064 0.000 58.216 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.064 0.000 58.216 0.152 ;
    END
  END O1[164]

  PIN I1[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.848 0.000 57.000 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.848 0.000 57.000 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.848 0.000 57.000 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.848 0.000 57.000 0.152 ;
    END
  END I1[164]

  PIN I1[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.544 0.000 56.696 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.544 0.000 56.696 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.544 0.000 56.696 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.544 0.000 56.696 0.152 ;
    END
  END I1[165]

  PIN I1[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.240 0.000 56.392 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.240 0.000 56.392 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.240 0.000 56.392 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.240 0.000 56.392 0.152 ;
    END
  END I1[166]

  PIN I1[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.936 0.000 56.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.936 0.000 56.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.936 0.000 56.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.936 0.000 56.088 0.152 ;
    END
  END I1[167]

  PIN O1[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.720 0.000 54.872 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.720 0.000 54.872 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.720 0.000 54.872 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.720 0.000 54.872 0.152 ;
    END
  END O1[171]

  PIN O1[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.416 0.000 54.568 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.416 0.000 54.568 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.416 0.000 54.568 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.416 0.000 54.568 0.152 ;
    END
  END O1[170]

  PIN O1[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.112 0.000 54.264 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.112 0.000 54.264 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.112 0.000 54.264 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.112 0.000 54.264 0.152 ;
    END
  END O1[169]

  PIN O1[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.808 0.000 53.960 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.808 0.000 53.960 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.808 0.000 53.960 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.808 0.000 53.960 0.152 ;
    END
  END O1[168]

  PIN I1[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.592 0.000 52.744 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.592 0.000 52.744 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.592 0.000 52.744 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.592 0.000 52.744 0.152 ;
    END
  END I1[168]

  PIN I1[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.288 0.000 52.440 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.288 0.000 52.440 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.288 0.000 52.440 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.288 0.000 52.440 0.152 ;
    END
  END I1[169]

  PIN I1[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.984 0.000 52.136 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.984 0.000 52.136 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.984 0.000 52.136 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.984 0.000 52.136 0.152 ;
    END
  END I1[170]

  PIN I1[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.680 0.000 51.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.680 0.000 51.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.680 0.000 51.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.680 0.000 51.832 0.152 ;
    END
  END I1[171]

  PIN O1[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
  END O1[175]

  PIN O1[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
  END O1[174]

  PIN O1[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
  END O1[173]

  PIN O1[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
  END O1[172]

  PIN I1[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.336 0.000 48.488 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.336 0.000 48.488 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.336 0.000 48.488 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.336 0.000 48.488 0.152 ;
    END
  END I1[172]

  PIN I1[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.032 0.000 48.184 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.032 0.000 48.184 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.032 0.000 48.184 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.032 0.000 48.184 0.152 ;
    END
  END I1[173]

  PIN I1[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.728 0.000 47.880 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.728 0.000 47.880 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.728 0.000 47.880 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.728 0.000 47.880 0.152 ;
    END
  END I1[174]

  PIN I1[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.424 0.000 47.576 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.424 0.000 47.576 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.424 0.000 47.576 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.424 0.000 47.576 0.152 ;
    END
  END I1[175]

  PIN O1[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
  END O1[179]

  PIN O1[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.904 0.000 46.056 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.904 0.000 46.056 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.904 0.000 46.056 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.904 0.000 46.056 0.152 ;
    END
  END O1[178]

  PIN O1[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.600 0.000 45.752 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.600 0.000 45.752 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.600 0.000 45.752 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.600 0.000 45.752 0.152 ;
    END
  END O1[177]

  PIN O1[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.296 0.000 45.448 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.296 0.000 45.448 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.296 0.000 45.448 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.296 0.000 45.448 0.152 ;
    END
  END O1[176]

  PIN I1[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
  END I1[176]

  PIN I1[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
  END I1[177]

  PIN I1[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
  END I1[178]

  PIN I1[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
  END I1[179]

  PIN O1[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.952 0.000 42.104 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.952 0.000 42.104 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.952 0.000 42.104 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.952 0.000 42.104 0.152 ;
    END
  END O1[183]

  PIN O1[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.648 0.000 41.800 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.648 0.000 41.800 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.648 0.000 41.800 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.648 0.000 41.800 0.152 ;
    END
  END O1[182]

  PIN O1[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.344 0.000 41.496 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.344 0.000 41.496 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.344 0.000 41.496 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.344 0.000 41.496 0.152 ;
    END
  END O1[181]

  PIN O1[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.040 0.000 41.192 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.040 0.000 41.192 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.040 0.000 41.192 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.040 0.000 41.192 0.152 ;
    END
  END O1[180]

  PIN I1[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.824 0.000 39.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.824 0.000 39.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.824 0.000 39.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.824 0.000 39.976 0.152 ;
    END
  END I1[180]

  PIN I1[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.520 0.000 39.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.520 0.000 39.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.520 0.000 39.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.520 0.000 39.672 0.152 ;
    END
  END I1[181]

  PIN I1[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
  END I1[182]

  PIN I1[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
  END I1[183]

  PIN O1[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
  END O1[187]

  PIN O1[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.392 0.000 37.544 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.392 0.000 37.544 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.392 0.000 37.544 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.392 0.000 37.544 0.152 ;
    END
  END O1[186]

  PIN O1[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
  END O1[185]

  PIN O1[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.784 0.000 36.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.784 0.000 36.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.784 0.000 36.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.784 0.000 36.936 0.152 ;
    END
  END O1[184]

  PIN I1[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.568 0.000 35.720 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.568 0.000 35.720 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.568 0.000 35.720 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.568 0.000 35.720 0.152 ;
    END
  END I1[184]

  PIN I1[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.264 0.000 35.416 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.264 0.000 35.416 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.264 0.000 35.416 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.264 0.000 35.416 0.152 ;
    END
  END I1[185]

  PIN I1[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
  END I1[186]

  PIN I1[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
  END I1[187]

  PIN O1[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.440 0.000 33.592 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.440 0.000 33.592 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.440 0.000 33.592 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.440 0.000 33.592 0.152 ;
    END
  END O1[191]

  PIN O1[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.136 0.000 33.288 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.136 0.000 33.288 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.136 0.000 33.288 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.136 0.000 33.288 0.152 ;
    END
  END O1[190]

  PIN O1[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.832 0.000 32.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.832 0.000 32.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.832 0.000 32.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.832 0.000 32.984 0.152 ;
    END
  END O1[189]

  PIN O1[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.528 0.000 32.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.528 0.000 32.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.528 0.000 32.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.528 0.000 32.680 0.152 ;
    END
  END O1[188]

  PIN I1[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.312 0.000 31.464 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.312 0.000 31.464 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.312 0.000 31.464 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.312 0.000 31.464 0.152 ;
    END
  END I1[188]

  PIN I1[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.008 0.000 31.160 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.008 0.000 31.160 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.008 0.000 31.160 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.008 0.000 31.160 0.152 ;
    END
  END I1[189]

  PIN I1[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.704 0.000 30.856 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.704 0.000 30.856 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.704 0.000 30.856 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.704 0.000 30.856 0.152 ;
    END
  END I1[190]

  PIN I1[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.400 0.000 30.552 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.400 0.000 30.552 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.400 0.000 30.552 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.400 0.000 30.552 0.152 ;
    END
  END I1[191]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 92.568 260.224 92.720 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 92.568 260.224 92.720 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 92.568 260.224 92.720 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 92.568 260.224 92.720 ;
    END
  END A1[0]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 88.920 260.224 89.072 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 88.920 260.224 89.072 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 88.920 260.224 89.072 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 88.920 260.224 89.072 ;
    END
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 85.272 260.224 85.424 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 85.272 260.224 85.424 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 85.272 260.224 85.424 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 85.272 260.224 85.424 ;
    END
  END A1[2]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 81.624 260.224 81.776 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 81.624 260.224 81.776 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 81.624 260.224 81.776 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 81.624 260.224 81.776 ;
    END
  END A1[3]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 77.976 260.224 78.128 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 77.976 260.224 78.128 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 77.976 260.224 78.128 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 77.976 260.224 78.128 ;
    END
  END A1[4]

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 74.328 260.224 74.480 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 74.328 260.224 74.480 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 74.328 260.224 74.480 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 74.328 260.224 74.480 ;
    END
  END A1[5]

  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 70.680 260.224 70.832 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 70.680 260.224 70.832 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 70.680 260.224 70.832 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 70.680 260.224 70.832 ;
    END
  END A1[6]

  PIN A1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 67.032 260.224 67.184 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 67.032 260.224 67.184 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 67.032 260.224 67.184 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 67.032 260.224 67.184 ;
    END
  END A1[7]

  PIN A1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 63.384 260.224 63.536 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 63.384 260.224 63.536 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 63.384 260.224 63.536 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 63.384 260.224 63.536 ;
    END
  END A1[8]

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 26.448 260.224 26.600 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 26.448 260.224 26.600 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 26.448 260.224 26.600 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 26.448 260.224 26.600 ;
    END
  END WEB1

  PIN WBM1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 25.232 260.224 25.384 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 25.232 260.224 25.384 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 25.232 260.224 25.384 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 25.232 260.224 25.384 ;
    END
  END WBM1[0]

  PIN WBM1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 24.016 260.224 24.168 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 24.016 260.224 24.168 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 24.016 260.224 24.168 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 24.016 260.224 24.168 ;
    END
  END WBM1[1]

  PIN WBM1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 22.800 260.224 22.952 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 22.800 260.224 22.952 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 22.800 260.224 22.952 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 22.800 260.224 22.952 ;
    END
  END WBM1[2]

  PIN WBM1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 21.584 260.224 21.736 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 21.584 260.224 21.736 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 21.584 260.224 21.736 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 21.584 260.224 21.736 ;
    END
  END WBM1[3]

  PIN WBM1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 20.368 260.224 20.520 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 20.368 260.224 20.520 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 20.368 260.224 20.520 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 20.368 260.224 20.520 ;
    END
  END WBM1[4]

  PIN WBM1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 19.152 260.224 19.304 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 19.152 260.224 19.304 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 19.152 260.224 19.304 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 19.152 260.224 19.304 ;
    END
  END WBM1[5]

  PIN WBM1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 17.936 260.224 18.088 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 17.936 260.224 18.088 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 17.936 260.224 18.088 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 17.936 260.224 18.088 ;
    END
  END WBM1[6]

  PIN WBM1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 16.720 260.224 16.872 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 16.720 260.224 16.872 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 16.720 260.224 16.872 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 16.720 260.224 16.872 ;
    END
  END WBM1[7]

  PIN WBM1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 15.504 260.224 15.656 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 15.504 260.224 15.656 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 15.504 260.224 15.656 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 15.504 260.224 15.656 ;
    END
  END WBM1[8]

  PIN WBM1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 14.288 260.224 14.440 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 14.288 260.224 14.440 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 14.288 260.224 14.440 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 14.288 260.224 14.440 ;
    END
  END WBM1[9]

  PIN WBM1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 13.072 260.224 13.224 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 13.072 260.224 13.224 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 13.072 260.224 13.224 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 13.072 260.224 13.224 ;
    END
  END WBM1[10]

  PIN WBM1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 11.856 260.224 12.008 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 11.856 260.224 12.008 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 11.856 260.224 12.008 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 11.856 260.224 12.008 ;
    END
  END WBM1[11]

  PIN WBM1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 10.640 260.224 10.792 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 10.640 260.224 10.792 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 10.640 260.224 10.792 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 10.640 260.224 10.792 ;
    END
  END WBM1[12]

  PIN WBM1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 9.424 260.224 9.576 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 9.424 260.224 9.576 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 9.424 260.224 9.576 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 9.424 260.224 9.576 ;
    END
  END WBM1[13]

  PIN WBM1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 8.208 260.224 8.360 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 8.208 260.224 8.360 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 8.208 260.224 8.360 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 8.208 260.224 8.360 ;
    END
  END WBM1[14]

  PIN WBM1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 6.992 260.224 7.144 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 6.992 260.224 7.144 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 6.992 260.224 7.144 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 6.992 260.224 7.144 ;
    END
  END WBM1[15]

  PIN WBM1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 5.776 260.224 5.928 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 5.776 260.224 5.928 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 5.776 260.224 5.928 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 5.776 260.224 5.928 ;
    END
  END WBM1[16]

  PIN WBM1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 4.560 260.224 4.712 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 4.560 260.224 4.712 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 4.560 260.224 4.712 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 4.560 260.224 4.712 ;
    END
  END WBM1[17]

  PIN WBM1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 3.344 260.224 3.496 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 3.344 260.224 3.496 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 3.344 260.224 3.496 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 3.344 260.224 3.496 ;
    END
  END WBM1[18]

  PIN WBM1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 2.128 260.224 2.280 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 2.128 260.224 2.280 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 2.128 260.224 2.280 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 2.128 260.224 2.280 ;
    END
  END WBM1[19]

  PIN WBM1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 0.912 260.224 1.064 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 0.912 260.224 1.064 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 0.912 260.224 1.064 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 0.912 260.224 1.064 ;
    END
  END WBM1[20]

  PIN WBM1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 -0.304 260.224 -0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 -0.304 260.224 -0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 -0.304 260.224 -0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 -0.304 260.224 -0.152 ;
    END
  END WBM1[21]

  PIN WBM1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 -1.520 260.224 -1.368 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 -1.520 260.224 -1.368 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 -1.520 260.224 -1.368 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 -1.520 260.224 -1.368 ;
    END
  END WBM1[22]

  PIN WBM1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 260.072 -2.736 260.224 -2.584 ;
    END
    PORT
      LAYER M3 ;
        RECT 260.072 -2.736 260.224 -2.584 ;
    END
    PORT
      LAYER M4 ;
        RECT 260.072 -2.736 260.224 -2.584 ;
    END
    PORT
      LAYER M5 ;
        RECT 260.072 -2.736 260.224 -2.584 ;
    END
  END WBM1[23]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 5.195 103.792 7.195 105.792 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.195 103.792 7.195 105.792 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.195 103.792 7.195 105.792 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M2 ;
        RECT 7.915 103.792 9.915 105.792 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.915 103.792 9.915 105.792 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.915 103.792 9.915 105.792 ;
    END
  END VSS

  OBS
    LAYER M2 ;
      RECT 237.424 0.000 260.224 0.304 ;
      RECT 236.208 0.000 236.968 0.304 ;
      RECT 234.992 0.000 235.752 0.304 ;
      RECT 233.776 0.000 234.536 0.304 ;
      RECT 231.648 0.000 232.408 0.304 ;
      RECT 229.520 0.000 230.280 0.304 ;
      RECT 227.392 0.000 228.152 0.304 ;
      RECT 225.264 0.000 226.024 0.304 ;
      RECT 223.136 0.000 223.896 0.304 ;
      RECT 221.008 0.000 221.768 0.304 ;
      RECT 218.880 0.000 219.640 0.304 ;
      RECT 216.752 0.000 217.512 0.304 ;
      RECT 214.624 0.000 215.384 0.304 ;
      RECT 212.496 0.000 213.256 0.304 ;
      RECT 210.368 0.000 211.128 0.304 ;
      RECT 208.240 0.000 209.000 0.304 ;
      RECT 206.112 0.000 206.872 0.304 ;
      RECT 203.984 0.000 204.744 0.304 ;
      RECT 201.856 0.000 202.616 0.304 ;
      RECT 199.728 0.000 200.488 0.304 ;
      RECT 197.600 0.000 198.360 0.304 ;
      RECT 195.472 0.000 196.232 0.304 ;
      RECT 193.344 0.000 194.104 0.304 ;
      RECT 191.216 0.000 191.976 0.304 ;
      RECT 189.088 0.000 189.848 0.304 ;
      RECT 186.960 0.000 187.720 0.304 ;
      RECT 184.832 0.000 185.592 0.304 ;
      RECT 182.704 0.000 183.464 0.304 ;
      RECT 180.576 0.000 181.336 0.304 ;
      RECT 178.448 0.000 179.208 0.304 ;
      RECT 176.320 0.000 177.080 0.304 ;
      RECT 174.192 0.000 174.952 0.304 ;
      RECT 172.064 0.000 172.824 0.304 ;
      RECT 169.936 0.000 170.696 0.304 ;
      RECT 167.808 0.000 168.568 0.304 ;
      RECT 165.680 0.000 166.440 0.304 ;
      RECT 163.552 0.000 164.312 0.304 ;
      RECT 161.424 0.000 162.184 0.304 ;
      RECT 159.296 0.000 160.056 0.304 ;
      RECT 157.168 0.000 157.928 0.304 ;
      RECT 155.040 0.000 155.800 0.304 ;
      RECT 152.912 0.000 153.672 0.304 ;
      RECT 150.784 0.000 151.544 0.304 ;
      RECT 148.656 0.000 149.416 0.304 ;
      RECT 146.528 0.000 147.288 0.304 ;
      RECT 144.400 0.000 145.160 0.304 ;
      RECT 142.272 0.000 143.032 0.304 ;
      RECT 140.144 0.000 140.904 0.304 ;
      RECT 138.016 0.000 138.776 0.304 ;
      RECT 135.888 0.000 136.648 0.304 ;
      RECT 133.760 0.000 134.520 0.304 ;
      RECT 131.632 0.000 132.392 0.304 ;
      RECT 129.504 0.000 130.264 0.304 ;
      RECT 127.376 0.000 128.136 0.304 ;
      RECT 125.248 0.000 126.008 0.304 ;
      RECT 123.120 0.000 123.880 0.304 ;
      RECT 120.992 0.000 121.752 0.304 ;
      RECT 118.864 0.000 119.624 0.304 ;
      RECT 116.736 0.000 117.496 0.304 ;
      RECT 114.608 0.000 115.368 0.304 ;
      RECT 112.480 0.000 113.240 0.304 ;
      RECT 110.352 0.000 111.112 0.304 ;
      RECT 108.224 0.000 108.984 0.304 ;
      RECT 106.096 0.000 106.856 0.304 ;
      RECT 103.968 0.000 104.728 0.304 ;
      RECT 101.840 0.000 102.600 0.304 ;
      RECT 99.712 0.000 100.472 0.304 ;
      RECT 97.584 0.000 98.344 0.304 ;
      RECT 95.456 0.000 96.216 0.304 ;
      RECT 93.328 0.000 94.088 0.304 ;
      RECT 91.200 0.000 91.960 0.304 ;
      RECT 89.072 0.000 89.832 0.304 ;
      RECT 86.944 0.000 87.704 0.304 ;
      RECT 84.816 0.000 85.576 0.304 ;
      RECT 82.688 0.000 83.448 0.304 ;
      RECT 80.560 0.000 81.320 0.304 ;
      RECT 78.432 0.000 79.192 0.304 ;
      RECT 76.304 0.000 77.064 0.304 ;
      RECT 74.176 0.000 74.936 0.304 ;
      RECT 72.048 0.000 72.808 0.304 ;
      RECT 69.920 0.000 70.680 0.304 ;
      RECT 67.792 0.000 68.552 0.304 ;
      RECT 65.664 0.000 66.424 0.304 ;
      RECT 63.536 0.000 64.296 0.304 ;
      RECT 61.408 0.000 62.168 0.304 ;
      RECT 59.280 0.000 60.040 0.304 ;
      RECT 57.152 0.000 57.912 0.304 ;
      RECT 55.024 0.000 55.784 0.304 ;
      RECT 52.896 0.000 53.656 0.304 ;
      RECT 50.768 0.000 51.528 0.304 ;
      RECT 48.640 0.000 49.400 0.304 ;
      RECT 46.512 0.000 47.272 0.304 ;
      RECT 44.384 0.000 45.144 0.304 ;
      RECT 42.256 0.000 43.016 0.304 ;
      RECT 40.128 0.000 40.888 0.304 ;
      RECT 38.000 0.000 38.760 0.304 ;
      RECT 35.872 0.000 36.632 0.304 ;
      RECT 33.744 0.000 34.504 0.304 ;
      RECT 31.616 0.000 32.376 0.304 ;
      RECT 0.000 0.000 30.248 0.304 ;
      RECT 259.920 92.872 260.224 103.640 ;
      RECT 259.920 89.224 260.224 92.416 ;
      RECT 259.920 85.576 260.224 88.768 ;
      RECT 259.920 81.928 260.224 85.120 ;
      RECT 259.920 78.280 260.224 81.472 ;
      RECT 259.920 74.632 260.224 77.824 ;
      RECT 259.920 70.984 260.224 74.176 ;
      RECT 259.920 67.336 260.224 70.528 ;
      RECT 259.920 63.688 260.224 66.880 ;
      RECT 259.920 26.752 260.224 63.232 ;
      RECT 259.920 25.536 260.224 26.296 ;
      RECT 259.920 24.320 260.224 25.080 ;
      RECT 259.920 23.104 260.224 23.864 ;
      RECT 259.920 21.888 260.224 22.648 ;
      RECT 259.920 20.672 260.224 21.432 ;
      RECT 259.920 19.456 260.224 20.216 ;
      RECT 259.920 18.240 260.224 19.000 ;
      RECT 259.920 17.024 260.224 17.784 ;
      RECT 259.920 15.808 260.224 16.568 ;
      RECT 259.920 14.592 260.224 15.352 ;
      RECT 259.920 13.376 260.224 14.136 ;
      RECT 259.920 12.160 260.224 12.920 ;
      RECT 259.920 10.944 260.224 11.704 ;
      RECT 259.920 9.728 260.224 10.488 ;
      RECT 259.920 8.512 260.224 9.272 ;
      RECT 259.920 7.296 260.224 8.056 ;
      RECT 259.920 6.080 260.224 6.840 ;
      RECT 259.920 4.864 260.224 5.624 ;
      RECT 259.920 3.648 260.224 4.408 ;
      RECT 259.920 2.432 260.224 3.192 ;
      RECT 259.920 1.216 260.224 1.976 ;
      RECT 259.920 -0.000 260.224 0.760 ;
      RECT 259.920 -1.216 260.224 -0.456 ;
      RECT 259.920 -2.432 260.224 -1.672 ;
      RECT 259.920 0.304 260.224 -2.888 ;
      RECT 0.000 103.640 5.043 105.792 ;
      RECT 7.355 103.640 7.763 105.792 ;
      RECT 10.067 103.640 260.224 105.792 ;
      RECT 0.000 0.304 259.920 103.640 ;
    LAYER M3 ;
      RECT 237.424 0.000 260.224 0.304 ;
      RECT 236.208 0.000 236.968 0.304 ;
      RECT 234.992 0.000 235.752 0.304 ;
      RECT 233.776 0.000 234.536 0.304 ;
      RECT 231.648 0.000 232.408 0.304 ;
      RECT 229.520 0.000 230.280 0.304 ;
      RECT 227.392 0.000 228.152 0.304 ;
      RECT 225.264 0.000 226.024 0.304 ;
      RECT 223.136 0.000 223.896 0.304 ;
      RECT 221.008 0.000 221.768 0.304 ;
      RECT 218.880 0.000 219.640 0.304 ;
      RECT 216.752 0.000 217.512 0.304 ;
      RECT 214.624 0.000 215.384 0.304 ;
      RECT 212.496 0.000 213.256 0.304 ;
      RECT 210.368 0.000 211.128 0.304 ;
      RECT 208.240 0.000 209.000 0.304 ;
      RECT 206.112 0.000 206.872 0.304 ;
      RECT 203.984 0.000 204.744 0.304 ;
      RECT 201.856 0.000 202.616 0.304 ;
      RECT 199.728 0.000 200.488 0.304 ;
      RECT 197.600 0.000 198.360 0.304 ;
      RECT 195.472 0.000 196.232 0.304 ;
      RECT 193.344 0.000 194.104 0.304 ;
      RECT 191.216 0.000 191.976 0.304 ;
      RECT 189.088 0.000 189.848 0.304 ;
      RECT 186.960 0.000 187.720 0.304 ;
      RECT 184.832 0.000 185.592 0.304 ;
      RECT 182.704 0.000 183.464 0.304 ;
      RECT 180.576 0.000 181.336 0.304 ;
      RECT 178.448 0.000 179.208 0.304 ;
      RECT 176.320 0.000 177.080 0.304 ;
      RECT 174.192 0.000 174.952 0.304 ;
      RECT 172.064 0.000 172.824 0.304 ;
      RECT 169.936 0.000 170.696 0.304 ;
      RECT 167.808 0.000 168.568 0.304 ;
      RECT 165.680 0.000 166.440 0.304 ;
      RECT 163.552 0.000 164.312 0.304 ;
      RECT 161.424 0.000 162.184 0.304 ;
      RECT 159.296 0.000 160.056 0.304 ;
      RECT 157.168 0.000 157.928 0.304 ;
      RECT 155.040 0.000 155.800 0.304 ;
      RECT 152.912 0.000 153.672 0.304 ;
      RECT 150.784 0.000 151.544 0.304 ;
      RECT 148.656 0.000 149.416 0.304 ;
      RECT 146.528 0.000 147.288 0.304 ;
      RECT 144.400 0.000 145.160 0.304 ;
      RECT 142.272 0.000 143.032 0.304 ;
      RECT 140.144 0.000 140.904 0.304 ;
      RECT 138.016 0.000 138.776 0.304 ;
      RECT 135.888 0.000 136.648 0.304 ;
      RECT 133.760 0.000 134.520 0.304 ;
      RECT 131.632 0.000 132.392 0.304 ;
      RECT 129.504 0.000 130.264 0.304 ;
      RECT 127.376 0.000 128.136 0.304 ;
      RECT 125.248 0.000 126.008 0.304 ;
      RECT 123.120 0.000 123.880 0.304 ;
      RECT 120.992 0.000 121.752 0.304 ;
      RECT 118.864 0.000 119.624 0.304 ;
      RECT 116.736 0.000 117.496 0.304 ;
      RECT 114.608 0.000 115.368 0.304 ;
      RECT 112.480 0.000 113.240 0.304 ;
      RECT 110.352 0.000 111.112 0.304 ;
      RECT 108.224 0.000 108.984 0.304 ;
      RECT 106.096 0.000 106.856 0.304 ;
      RECT 103.968 0.000 104.728 0.304 ;
      RECT 101.840 0.000 102.600 0.304 ;
      RECT 99.712 0.000 100.472 0.304 ;
      RECT 97.584 0.000 98.344 0.304 ;
      RECT 95.456 0.000 96.216 0.304 ;
      RECT 93.328 0.000 94.088 0.304 ;
      RECT 91.200 0.000 91.960 0.304 ;
      RECT 89.072 0.000 89.832 0.304 ;
      RECT 86.944 0.000 87.704 0.304 ;
      RECT 84.816 0.000 85.576 0.304 ;
      RECT 82.688 0.000 83.448 0.304 ;
      RECT 80.560 0.000 81.320 0.304 ;
      RECT 78.432 0.000 79.192 0.304 ;
      RECT 76.304 0.000 77.064 0.304 ;
      RECT 74.176 0.000 74.936 0.304 ;
      RECT 72.048 0.000 72.808 0.304 ;
      RECT 69.920 0.000 70.680 0.304 ;
      RECT 67.792 0.000 68.552 0.304 ;
      RECT 65.664 0.000 66.424 0.304 ;
      RECT 63.536 0.000 64.296 0.304 ;
      RECT 61.408 0.000 62.168 0.304 ;
      RECT 59.280 0.000 60.040 0.304 ;
      RECT 57.152 0.000 57.912 0.304 ;
      RECT 55.024 0.000 55.784 0.304 ;
      RECT 52.896 0.000 53.656 0.304 ;
      RECT 50.768 0.000 51.528 0.304 ;
      RECT 48.640 0.000 49.400 0.304 ;
      RECT 46.512 0.000 47.272 0.304 ;
      RECT 44.384 0.000 45.144 0.304 ;
      RECT 42.256 0.000 43.016 0.304 ;
      RECT 40.128 0.000 40.888 0.304 ;
      RECT 38.000 0.000 38.760 0.304 ;
      RECT 35.872 0.000 36.632 0.304 ;
      RECT 33.744 0.000 34.504 0.304 ;
      RECT 31.616 0.000 32.376 0.304 ;
      RECT 0.000 0.000 30.248 0.304 ;
      RECT 259.920 92.872 260.224 103.640 ;
      RECT 259.920 89.224 260.224 92.416 ;
      RECT 259.920 85.576 260.224 88.768 ;
      RECT 259.920 81.928 260.224 85.120 ;
      RECT 259.920 78.280 260.224 81.472 ;
      RECT 259.920 74.632 260.224 77.824 ;
      RECT 259.920 70.984 260.224 74.176 ;
      RECT 259.920 67.336 260.224 70.528 ;
      RECT 259.920 63.688 260.224 66.880 ;
      RECT 259.920 26.752 260.224 63.232 ;
      RECT 259.920 25.536 260.224 26.296 ;
      RECT 259.920 24.320 260.224 25.080 ;
      RECT 259.920 23.104 260.224 23.864 ;
      RECT 259.920 21.888 260.224 22.648 ;
      RECT 259.920 20.672 260.224 21.432 ;
      RECT 259.920 19.456 260.224 20.216 ;
      RECT 259.920 18.240 260.224 19.000 ;
      RECT 259.920 17.024 260.224 17.784 ;
      RECT 259.920 15.808 260.224 16.568 ;
      RECT 259.920 14.592 260.224 15.352 ;
      RECT 259.920 13.376 260.224 14.136 ;
      RECT 259.920 12.160 260.224 12.920 ;
      RECT 259.920 10.944 260.224 11.704 ;
      RECT 259.920 9.728 260.224 10.488 ;
      RECT 259.920 8.512 260.224 9.272 ;
      RECT 259.920 7.296 260.224 8.056 ;
      RECT 259.920 6.080 260.224 6.840 ;
      RECT 259.920 4.864 260.224 5.624 ;
      RECT 259.920 3.648 260.224 4.408 ;
      RECT 259.920 2.432 260.224 3.192 ;
      RECT 259.920 1.216 260.224 1.976 ;
      RECT 259.920 -0.000 260.224 0.760 ;
      RECT 259.920 -1.216 260.224 -0.456 ;
      RECT 259.920 -2.432 260.224 -1.672 ;
      RECT 259.920 0.304 260.224 -2.888 ;
      RECT 0.000 103.640 5.043 105.792 ;
      RECT 7.355 103.640 7.763 105.792 ;
      RECT 10.067 103.640 260.224 105.792 ;
      RECT 0.000 0.304 259.920 103.640 ;
    LAYER M4 ;
      RECT 237.424 0.000 260.224 0.304 ;
      RECT 236.208 0.000 236.968 0.304 ;
      RECT 234.992 0.000 235.752 0.304 ;
      RECT 233.776 0.000 234.536 0.304 ;
      RECT 231.648 0.000 232.408 0.304 ;
      RECT 229.520 0.000 230.280 0.304 ;
      RECT 227.392 0.000 228.152 0.304 ;
      RECT 225.264 0.000 226.024 0.304 ;
      RECT 223.136 0.000 223.896 0.304 ;
      RECT 221.008 0.000 221.768 0.304 ;
      RECT 218.880 0.000 219.640 0.304 ;
      RECT 216.752 0.000 217.512 0.304 ;
      RECT 214.624 0.000 215.384 0.304 ;
      RECT 212.496 0.000 213.256 0.304 ;
      RECT 210.368 0.000 211.128 0.304 ;
      RECT 208.240 0.000 209.000 0.304 ;
      RECT 206.112 0.000 206.872 0.304 ;
      RECT 203.984 0.000 204.744 0.304 ;
      RECT 201.856 0.000 202.616 0.304 ;
      RECT 199.728 0.000 200.488 0.304 ;
      RECT 197.600 0.000 198.360 0.304 ;
      RECT 195.472 0.000 196.232 0.304 ;
      RECT 193.344 0.000 194.104 0.304 ;
      RECT 191.216 0.000 191.976 0.304 ;
      RECT 189.088 0.000 189.848 0.304 ;
      RECT 186.960 0.000 187.720 0.304 ;
      RECT 184.832 0.000 185.592 0.304 ;
      RECT 182.704 0.000 183.464 0.304 ;
      RECT 180.576 0.000 181.336 0.304 ;
      RECT 178.448 0.000 179.208 0.304 ;
      RECT 176.320 0.000 177.080 0.304 ;
      RECT 174.192 0.000 174.952 0.304 ;
      RECT 172.064 0.000 172.824 0.304 ;
      RECT 169.936 0.000 170.696 0.304 ;
      RECT 167.808 0.000 168.568 0.304 ;
      RECT 165.680 0.000 166.440 0.304 ;
      RECT 163.552 0.000 164.312 0.304 ;
      RECT 161.424 0.000 162.184 0.304 ;
      RECT 159.296 0.000 160.056 0.304 ;
      RECT 157.168 0.000 157.928 0.304 ;
      RECT 155.040 0.000 155.800 0.304 ;
      RECT 152.912 0.000 153.672 0.304 ;
      RECT 150.784 0.000 151.544 0.304 ;
      RECT 148.656 0.000 149.416 0.304 ;
      RECT 146.528 0.000 147.288 0.304 ;
      RECT 144.400 0.000 145.160 0.304 ;
      RECT 142.272 0.000 143.032 0.304 ;
      RECT 140.144 0.000 140.904 0.304 ;
      RECT 138.016 0.000 138.776 0.304 ;
      RECT 135.888 0.000 136.648 0.304 ;
      RECT 133.760 0.000 134.520 0.304 ;
      RECT 131.632 0.000 132.392 0.304 ;
      RECT 129.504 0.000 130.264 0.304 ;
      RECT 127.376 0.000 128.136 0.304 ;
      RECT 125.248 0.000 126.008 0.304 ;
      RECT 123.120 0.000 123.880 0.304 ;
      RECT 120.992 0.000 121.752 0.304 ;
      RECT 118.864 0.000 119.624 0.304 ;
      RECT 116.736 0.000 117.496 0.304 ;
      RECT 114.608 0.000 115.368 0.304 ;
      RECT 112.480 0.000 113.240 0.304 ;
      RECT 110.352 0.000 111.112 0.304 ;
      RECT 108.224 0.000 108.984 0.304 ;
      RECT 106.096 0.000 106.856 0.304 ;
      RECT 103.968 0.000 104.728 0.304 ;
      RECT 101.840 0.000 102.600 0.304 ;
      RECT 99.712 0.000 100.472 0.304 ;
      RECT 97.584 0.000 98.344 0.304 ;
      RECT 95.456 0.000 96.216 0.304 ;
      RECT 93.328 0.000 94.088 0.304 ;
      RECT 91.200 0.000 91.960 0.304 ;
      RECT 89.072 0.000 89.832 0.304 ;
      RECT 86.944 0.000 87.704 0.304 ;
      RECT 84.816 0.000 85.576 0.304 ;
      RECT 82.688 0.000 83.448 0.304 ;
      RECT 80.560 0.000 81.320 0.304 ;
      RECT 78.432 0.000 79.192 0.304 ;
      RECT 76.304 0.000 77.064 0.304 ;
      RECT 74.176 0.000 74.936 0.304 ;
      RECT 72.048 0.000 72.808 0.304 ;
      RECT 69.920 0.000 70.680 0.304 ;
      RECT 67.792 0.000 68.552 0.304 ;
      RECT 65.664 0.000 66.424 0.304 ;
      RECT 63.536 0.000 64.296 0.304 ;
      RECT 61.408 0.000 62.168 0.304 ;
      RECT 59.280 0.000 60.040 0.304 ;
      RECT 57.152 0.000 57.912 0.304 ;
      RECT 55.024 0.000 55.784 0.304 ;
      RECT 52.896 0.000 53.656 0.304 ;
      RECT 50.768 0.000 51.528 0.304 ;
      RECT 48.640 0.000 49.400 0.304 ;
      RECT 46.512 0.000 47.272 0.304 ;
      RECT 44.384 0.000 45.144 0.304 ;
      RECT 42.256 0.000 43.016 0.304 ;
      RECT 40.128 0.000 40.888 0.304 ;
      RECT 38.000 0.000 38.760 0.304 ;
      RECT 35.872 0.000 36.632 0.304 ;
      RECT 33.744 0.000 34.504 0.304 ;
      RECT 31.616 0.000 32.376 0.304 ;
      RECT 0.000 0.000 30.248 0.304 ;
      RECT 259.920 92.872 260.224 103.640 ;
      RECT 259.920 89.224 260.224 92.416 ;
      RECT 259.920 85.576 260.224 88.768 ;
      RECT 259.920 81.928 260.224 85.120 ;
      RECT 259.920 78.280 260.224 81.472 ;
      RECT 259.920 74.632 260.224 77.824 ;
      RECT 259.920 70.984 260.224 74.176 ;
      RECT 259.920 67.336 260.224 70.528 ;
      RECT 259.920 63.688 260.224 66.880 ;
      RECT 259.920 26.752 260.224 63.232 ;
      RECT 259.920 25.536 260.224 26.296 ;
      RECT 259.920 24.320 260.224 25.080 ;
      RECT 259.920 23.104 260.224 23.864 ;
      RECT 259.920 21.888 260.224 22.648 ;
      RECT 259.920 20.672 260.224 21.432 ;
      RECT 259.920 19.456 260.224 20.216 ;
      RECT 259.920 18.240 260.224 19.000 ;
      RECT 259.920 17.024 260.224 17.784 ;
      RECT 259.920 15.808 260.224 16.568 ;
      RECT 259.920 14.592 260.224 15.352 ;
      RECT 259.920 13.376 260.224 14.136 ;
      RECT 259.920 12.160 260.224 12.920 ;
      RECT 259.920 10.944 260.224 11.704 ;
      RECT 259.920 9.728 260.224 10.488 ;
      RECT 259.920 8.512 260.224 9.272 ;
      RECT 259.920 7.296 260.224 8.056 ;
      RECT 259.920 6.080 260.224 6.840 ;
      RECT 259.920 4.864 260.224 5.624 ;
      RECT 259.920 3.648 260.224 4.408 ;
      RECT 259.920 2.432 260.224 3.192 ;
      RECT 259.920 1.216 260.224 1.976 ;
      RECT 259.920 -0.000 260.224 0.760 ;
      RECT 259.920 -1.216 260.224 -0.456 ;
      RECT 259.920 -2.432 260.224 -1.672 ;
      RECT 259.920 0.304 260.224 -2.888 ;
      RECT 0.000 103.640 5.043 105.792 ;
      RECT 7.355 103.640 7.763 105.792 ;
      RECT 10.067 103.640 260.224 105.792 ;
      RECT 0.000 0.304 259.920 103.640 ;
    LAYER M5 ;
      RECT 237.424 0.000 260.224 0.304 ;
      RECT 236.208 0.000 236.968 0.304 ;
      RECT 234.992 0.000 235.752 0.304 ;
      RECT 233.776 0.000 234.536 0.304 ;
      RECT 231.648 0.000 232.408 0.304 ;
      RECT 229.520 0.000 230.280 0.304 ;
      RECT 227.392 0.000 228.152 0.304 ;
      RECT 225.264 0.000 226.024 0.304 ;
      RECT 223.136 0.000 223.896 0.304 ;
      RECT 221.008 0.000 221.768 0.304 ;
      RECT 218.880 0.000 219.640 0.304 ;
      RECT 216.752 0.000 217.512 0.304 ;
      RECT 214.624 0.000 215.384 0.304 ;
      RECT 212.496 0.000 213.256 0.304 ;
      RECT 210.368 0.000 211.128 0.304 ;
      RECT 208.240 0.000 209.000 0.304 ;
      RECT 206.112 0.000 206.872 0.304 ;
      RECT 203.984 0.000 204.744 0.304 ;
      RECT 201.856 0.000 202.616 0.304 ;
      RECT 199.728 0.000 200.488 0.304 ;
      RECT 197.600 0.000 198.360 0.304 ;
      RECT 195.472 0.000 196.232 0.304 ;
      RECT 193.344 0.000 194.104 0.304 ;
      RECT 191.216 0.000 191.976 0.304 ;
      RECT 189.088 0.000 189.848 0.304 ;
      RECT 186.960 0.000 187.720 0.304 ;
      RECT 184.832 0.000 185.592 0.304 ;
      RECT 182.704 0.000 183.464 0.304 ;
      RECT 180.576 0.000 181.336 0.304 ;
      RECT 178.448 0.000 179.208 0.304 ;
      RECT 176.320 0.000 177.080 0.304 ;
      RECT 174.192 0.000 174.952 0.304 ;
      RECT 172.064 0.000 172.824 0.304 ;
      RECT 169.936 0.000 170.696 0.304 ;
      RECT 167.808 0.000 168.568 0.304 ;
      RECT 165.680 0.000 166.440 0.304 ;
      RECT 163.552 0.000 164.312 0.304 ;
      RECT 161.424 0.000 162.184 0.304 ;
      RECT 159.296 0.000 160.056 0.304 ;
      RECT 157.168 0.000 157.928 0.304 ;
      RECT 155.040 0.000 155.800 0.304 ;
      RECT 152.912 0.000 153.672 0.304 ;
      RECT 150.784 0.000 151.544 0.304 ;
      RECT 148.656 0.000 149.416 0.304 ;
      RECT 146.528 0.000 147.288 0.304 ;
      RECT 144.400 0.000 145.160 0.304 ;
      RECT 142.272 0.000 143.032 0.304 ;
      RECT 140.144 0.000 140.904 0.304 ;
      RECT 138.016 0.000 138.776 0.304 ;
      RECT 135.888 0.000 136.648 0.304 ;
      RECT 133.760 0.000 134.520 0.304 ;
      RECT 131.632 0.000 132.392 0.304 ;
      RECT 129.504 0.000 130.264 0.304 ;
      RECT 127.376 0.000 128.136 0.304 ;
      RECT 125.248 0.000 126.008 0.304 ;
      RECT 123.120 0.000 123.880 0.304 ;
      RECT 120.992 0.000 121.752 0.304 ;
      RECT 118.864 0.000 119.624 0.304 ;
      RECT 116.736 0.000 117.496 0.304 ;
      RECT 114.608 0.000 115.368 0.304 ;
      RECT 112.480 0.000 113.240 0.304 ;
      RECT 110.352 0.000 111.112 0.304 ;
      RECT 108.224 0.000 108.984 0.304 ;
      RECT 106.096 0.000 106.856 0.304 ;
      RECT 103.968 0.000 104.728 0.304 ;
      RECT 101.840 0.000 102.600 0.304 ;
      RECT 99.712 0.000 100.472 0.304 ;
      RECT 97.584 0.000 98.344 0.304 ;
      RECT 95.456 0.000 96.216 0.304 ;
      RECT 93.328 0.000 94.088 0.304 ;
      RECT 91.200 0.000 91.960 0.304 ;
      RECT 89.072 0.000 89.832 0.304 ;
      RECT 86.944 0.000 87.704 0.304 ;
      RECT 84.816 0.000 85.576 0.304 ;
      RECT 82.688 0.000 83.448 0.304 ;
      RECT 80.560 0.000 81.320 0.304 ;
      RECT 78.432 0.000 79.192 0.304 ;
      RECT 76.304 0.000 77.064 0.304 ;
      RECT 74.176 0.000 74.936 0.304 ;
      RECT 72.048 0.000 72.808 0.304 ;
      RECT 69.920 0.000 70.680 0.304 ;
      RECT 67.792 0.000 68.552 0.304 ;
      RECT 65.664 0.000 66.424 0.304 ;
      RECT 63.536 0.000 64.296 0.304 ;
      RECT 61.408 0.000 62.168 0.304 ;
      RECT 59.280 0.000 60.040 0.304 ;
      RECT 57.152 0.000 57.912 0.304 ;
      RECT 55.024 0.000 55.784 0.304 ;
      RECT 52.896 0.000 53.656 0.304 ;
      RECT 50.768 0.000 51.528 0.304 ;
      RECT 48.640 0.000 49.400 0.304 ;
      RECT 46.512 0.000 47.272 0.304 ;
      RECT 44.384 0.000 45.144 0.304 ;
      RECT 42.256 0.000 43.016 0.304 ;
      RECT 40.128 0.000 40.888 0.304 ;
      RECT 38.000 0.000 38.760 0.304 ;
      RECT 35.872 0.000 36.632 0.304 ;
      RECT 33.744 0.000 34.504 0.304 ;
      RECT 31.616 0.000 32.376 0.304 ;
      RECT 0.000 0.000 30.248 0.304 ;
      RECT 259.920 92.872 260.224 103.640 ;
      RECT 259.920 89.224 260.224 92.416 ;
      RECT 259.920 85.576 260.224 88.768 ;
      RECT 259.920 81.928 260.224 85.120 ;
      RECT 259.920 78.280 260.224 81.472 ;
      RECT 259.920 74.632 260.224 77.824 ;
      RECT 259.920 70.984 260.224 74.176 ;
      RECT 259.920 67.336 260.224 70.528 ;
      RECT 259.920 63.688 260.224 66.880 ;
      RECT 259.920 26.752 260.224 63.232 ;
      RECT 259.920 25.536 260.224 26.296 ;
      RECT 259.920 24.320 260.224 25.080 ;
      RECT 259.920 23.104 260.224 23.864 ;
      RECT 259.920 21.888 260.224 22.648 ;
      RECT 259.920 20.672 260.224 21.432 ;
      RECT 259.920 19.456 260.224 20.216 ;
      RECT 259.920 18.240 260.224 19.000 ;
      RECT 259.920 17.024 260.224 17.784 ;
      RECT 259.920 15.808 260.224 16.568 ;
      RECT 259.920 14.592 260.224 15.352 ;
      RECT 259.920 13.376 260.224 14.136 ;
      RECT 259.920 12.160 260.224 12.920 ;
      RECT 259.920 10.944 260.224 11.704 ;
      RECT 259.920 9.728 260.224 10.488 ;
      RECT 259.920 8.512 260.224 9.272 ;
      RECT 259.920 7.296 260.224 8.056 ;
      RECT 259.920 6.080 260.224 6.840 ;
      RECT 259.920 4.864 260.224 5.624 ;
      RECT 259.920 3.648 260.224 4.408 ;
      RECT 259.920 2.432 260.224 3.192 ;
      RECT 259.920 1.216 260.224 1.976 ;
      RECT 259.920 -0.000 260.224 0.760 ;
      RECT 259.920 -1.216 260.224 -0.456 ;
      RECT 259.920 -2.432 260.224 -1.672 ;
      RECT 259.920 0.304 260.224 -2.888 ;
      RECT 0.000 103.640 5.043 105.792 ;
      RECT 7.355 103.640 7.763 105.792 ;
      RECT 10.067 103.640 260.224 105.792 ;
      RECT 0.000 0.304 259.920 103.640 ;
  END

END sram6t512x192

END LIBRARY
