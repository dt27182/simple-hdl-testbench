VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram6t128x48
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 68.096 BY 38.912 ;
  SYMMETRY X Y R90 ;

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.016 0.000 62.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.016 0.000 62.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.016 0.000 62.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.016 0.000 62.168 0.152 ;
    END
  END CE1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.800 0.000 60.952 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.800 0.000 60.952 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.800 0.000 60.952 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.800 0.000 60.952 0.152 ;
    END
  END CSB1

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.584 0.000 59.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.584 0.000 59.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.584 0.000 59.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.584 0.000 59.736 0.152 ;
    END
  END OEB1

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.368 0.000 58.520 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.368 0.000 58.520 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.368 0.000 58.520 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.368 0.000 58.520 0.152 ;
    END
  END O1[3]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.064 0.000 58.216 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.064 0.000 58.216 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.064 0.000 58.216 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.064 0.000 58.216 0.152 ;
    END
  END O1[2]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.760 0.000 57.912 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.760 0.000 57.912 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.760 0.000 57.912 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.760 0.000 57.912 0.152 ;
    END
  END O1[1]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.456 0.000 57.608 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.456 0.000 57.608 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.456 0.000 57.608 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.456 0.000 57.608 0.152 ;
    END
  END O1[0]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.240 0.000 56.392 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.240 0.000 56.392 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.240 0.000 56.392 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.240 0.000 56.392 0.152 ;
    END
  END I1[0]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.936 0.000 56.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.936 0.000 56.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.936 0.000 56.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.936 0.000 56.088 0.152 ;
    END
  END I1[1]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.632 0.000 55.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.632 0.000 55.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.632 0.000 55.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.632 0.000 55.784 0.152 ;
    END
  END I1[2]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.328 0.000 55.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.328 0.000 55.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.328 0.000 55.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.328 0.000 55.480 0.152 ;
    END
  END I1[3]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.112 0.000 54.264 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.112 0.000 54.264 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.112 0.000 54.264 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.112 0.000 54.264 0.152 ;
    END
  END O1[7]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.808 0.000 53.960 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.808 0.000 53.960 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.808 0.000 53.960 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.808 0.000 53.960 0.152 ;
    END
  END O1[6]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.504 0.000 53.656 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.504 0.000 53.656 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.504 0.000 53.656 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.504 0.000 53.656 0.152 ;
    END
  END O1[5]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.200 0.000 53.352 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.200 0.000 53.352 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.200 0.000 53.352 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.200 0.000 53.352 0.152 ;
    END
  END O1[4]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.984 0.000 52.136 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.984 0.000 52.136 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.984 0.000 52.136 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.984 0.000 52.136 0.152 ;
    END
  END I1[4]

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.680 0.000 51.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.680 0.000 51.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.680 0.000 51.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.680 0.000 51.832 0.152 ;
    END
  END I1[5]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
  END I1[6]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
  END I1[7]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
  END O1[11]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
  END O1[10]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
  END O1[9]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.944 0.000 49.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.944 0.000 49.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.944 0.000 49.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.944 0.000 49.096 0.152 ;
    END
  END O1[8]

  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.728 0.000 47.880 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.728 0.000 47.880 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.728 0.000 47.880 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.728 0.000 47.880 0.152 ;
    END
  END I1[8]

  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.424 0.000 47.576 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.424 0.000 47.576 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.424 0.000 47.576 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.424 0.000 47.576 0.152 ;
    END
  END I1[9]

  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
  END I1[10]

  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
  END I1[11]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.600 0.000 45.752 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.600 0.000 45.752 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.600 0.000 45.752 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.600 0.000 45.752 0.152 ;
    END
  END O1[15]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.296 0.000 45.448 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.296 0.000 45.448 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.296 0.000 45.448 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.296 0.000 45.448 0.152 ;
    END
  END O1[14]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.992 0.000 45.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.992 0.000 45.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.992 0.000 45.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.992 0.000 45.144 0.152 ;
    END
  END O1[13]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
  END O1[12]

  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
  END I1[12]

  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
  END I1[13]

  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.864 0.000 43.016 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.864 0.000 43.016 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.864 0.000 43.016 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.864 0.000 43.016 0.152 ;
    END
  END I1[14]

  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.560 0.000 42.712 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.560 0.000 42.712 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.560 0.000 42.712 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.560 0.000 42.712 0.152 ;
    END
  END I1[15]

  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.344 0.000 41.496 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.344 0.000 41.496 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.344 0.000 41.496 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.344 0.000 41.496 0.152 ;
    END
  END O1[19]

  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.040 0.000 41.192 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.040 0.000 41.192 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.040 0.000 41.192 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.040 0.000 41.192 0.152 ;
    END
  END O1[18]

  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.736 0.000 40.888 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.736 0.000 40.888 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.736 0.000 40.888 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.736 0.000 40.888 0.152 ;
    END
  END O1[17]

  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.432 0.000 40.584 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.432 0.000 40.584 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.432 0.000 40.584 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.432 0.000 40.584 0.152 ;
    END
  END O1[16]

  PIN I1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
  END I1[16]

  PIN I1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
  END I1[17]

  PIN I1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
  END I1[18]

  PIN I1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
  END I1[19]

  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.088 0.000 37.240 0.152 ;
    END
  END O1[23]

  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.784 0.000 36.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.784 0.000 36.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.784 0.000 36.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.784 0.000 36.936 0.152 ;
    END
  END O1[22]

  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.480 0.000 36.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.480 0.000 36.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.480 0.000 36.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.480 0.000 36.632 0.152 ;
    END
  END O1[21]

  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.176 0.000 36.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.176 0.000 36.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.176 0.000 36.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.176 0.000 36.328 0.152 ;
    END
  END O1[20]

  PIN I1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
  END I1[20]

  PIN I1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
  END I1[21]

  PIN I1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
  END I1[22]

  PIN I1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
  END I1[23]

  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.832 0.000 32.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.832 0.000 32.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.832 0.000 32.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.832 0.000 32.984 0.152 ;
    END
  END O1[27]

  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.528 0.000 32.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.528 0.000 32.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.528 0.000 32.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.528 0.000 32.680 0.152 ;
    END
  END O1[26]

  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.224 0.000 32.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.224 0.000 32.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.224 0.000 32.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.224 0.000 32.376 0.152 ;
    END
  END O1[25]

  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
  END O1[24]

  PIN I1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.704 0.000 30.856 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.704 0.000 30.856 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.704 0.000 30.856 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.704 0.000 30.856 0.152 ;
    END
  END I1[24]

  PIN I1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.400 0.000 30.552 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.400 0.000 30.552 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.400 0.000 30.552 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.400 0.000 30.552 0.152 ;
    END
  END I1[25]

  PIN I1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.096 0.000 30.248 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.096 0.000 30.248 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.096 0.000 30.248 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.096 0.000 30.248 0.152 ;
    END
  END I1[26]

  PIN I1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.792 0.000 29.944 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.792 0.000 29.944 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.792 0.000 29.944 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.792 0.000 29.944 0.152 ;
    END
  END I1[27]

  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.576 0.000 28.728 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.576 0.000 28.728 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.576 0.000 28.728 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.576 0.000 28.728 0.152 ;
    END
  END O1[31]

  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.272 0.000 28.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.272 0.000 28.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.272 0.000 28.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.272 0.000 28.424 0.152 ;
    END
  END O1[30]

  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
  END O1[29]

  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.664 0.000 27.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.664 0.000 27.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.664 0.000 27.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.664 0.000 27.816 0.152 ;
    END
  END O1[28]

  PIN I1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.448 0.000 26.600 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.448 0.000 26.600 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.448 0.000 26.600 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.448 0.000 26.600 0.152 ;
    END
  END I1[28]

  PIN I1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.144 0.000 26.296 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.144 0.000 26.296 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.144 0.000 26.296 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.144 0.000 26.296 0.152 ;
    END
  END I1[29]

  PIN I1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.840 0.000 25.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.840 0.000 25.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.840 0.000 25.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.840 0.000 25.992 0.152 ;
    END
  END I1[30]

  PIN I1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.536 0.000 25.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.536 0.000 25.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.536 0.000 25.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.536 0.000 25.688 0.152 ;
    END
  END I1[31]

  PIN O1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.320 0.000 24.472 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.320 0.000 24.472 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.320 0.000 24.472 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.320 0.000 24.472 0.152 ;
    END
  END O1[35]

  PIN O1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.016 0.000 24.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.016 0.000 24.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.016 0.000 24.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.016 0.000 24.168 0.152 ;
    END
  END O1[34]

  PIN O1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.712 0.000 23.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.712 0.000 23.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.712 0.000 23.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.712 0.000 23.864 0.152 ;
    END
  END O1[33]

  PIN O1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.408 0.000 23.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.408 0.000 23.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.408 0.000 23.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.408 0.000 23.560 0.152 ;
    END
  END O1[32]

  PIN I1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.192 0.000 22.344 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.192 0.000 22.344 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.192 0.000 22.344 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.192 0.000 22.344 0.152 ;
    END
  END I1[32]

  PIN I1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.888 0.000 22.040 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.888 0.000 22.040 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.888 0.000 22.040 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.888 0.000 22.040 0.152 ;
    END
  END I1[33]

  PIN I1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.584 0.000 21.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.584 0.000 21.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.584 0.000 21.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.584 0.000 21.736 0.152 ;
    END
  END I1[34]

  PIN I1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.280 0.000 21.432 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.280 0.000 21.432 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.280 0.000 21.432 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.280 0.000 21.432 0.152 ;
    END
  END I1[35]

  PIN O1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.064 0.000 20.216 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.064 0.000 20.216 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.064 0.000 20.216 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.064 0.000 20.216 0.152 ;
    END
  END O1[39]

  PIN O1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.760 0.000 19.912 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.760 0.000 19.912 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.760 0.000 19.912 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.760 0.000 19.912 0.152 ;
    END
  END O1[38]

  PIN O1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.456 0.000 19.608 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.456 0.000 19.608 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.456 0.000 19.608 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.456 0.000 19.608 0.152 ;
    END
  END O1[37]

  PIN O1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.152 0.000 19.304 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.152 0.000 19.304 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.152 0.000 19.304 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.152 0.000 19.304 0.152 ;
    END
  END O1[36]

  PIN I1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.936 0.000 18.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.936 0.000 18.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.936 0.000 18.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.936 0.000 18.088 0.152 ;
    END
  END I1[36]

  PIN I1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.632 0.000 17.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.632 0.000 17.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.632 0.000 17.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.632 0.000 17.784 0.152 ;
    END
  END I1[37]

  PIN I1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.328 0.000 17.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.328 0.000 17.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.328 0.000 17.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.328 0.000 17.480 0.152 ;
    END
  END I1[38]

  PIN I1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.024 0.000 17.176 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.024 0.000 17.176 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.024 0.000 17.176 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.024 0.000 17.176 0.152 ;
    END
  END I1[39]

  PIN O1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.808 0.000 15.960 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.808 0.000 15.960 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.808 0.000 15.960 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.808 0.000 15.960 0.152 ;
    END
  END O1[43]

  PIN O1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.504 0.000 15.656 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.504 0.000 15.656 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.504 0.000 15.656 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.504 0.000 15.656 0.152 ;
    END
  END O1[42]

  PIN O1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.200 0.000 15.352 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.200 0.000 15.352 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.200 0.000 15.352 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.200 0.000 15.352 0.152 ;
    END
  END O1[41]

  PIN O1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.896 0.000 15.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 14.896 0.000 15.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 14.896 0.000 15.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.896 0.000 15.048 0.152 ;
    END
  END O1[40]

  PIN I1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.680 0.000 13.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.680 0.000 13.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.680 0.000 13.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.680 0.000 13.832 0.152 ;
    END
  END I1[40]

  PIN I1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.376 0.000 13.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.376 0.000 13.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.376 0.000 13.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.376 0.000 13.528 0.152 ;
    END
  END I1[41]

  PIN I1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.072 0.000 13.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.072 0.000 13.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.072 0.000 13.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.072 0.000 13.224 0.152 ;
    END
  END I1[42]

  PIN I1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.768 0.000 12.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.768 0.000 12.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.768 0.000 12.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.768 0.000 12.920 0.152 ;
    END
  END I1[43]

  PIN O1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.552 0.000 11.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.552 0.000 11.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.552 0.000 11.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.552 0.000 11.704 0.152 ;
    END
  END O1[47]

  PIN O1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.248 0.000 11.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.248 0.000 11.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.248 0.000 11.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.248 0.000 11.400 0.152 ;
    END
  END O1[46]

  PIN O1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.944 0.000 11.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.944 0.000 11.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.944 0.000 11.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.944 0.000 11.096 0.152 ;
    END
  END O1[45]

  PIN O1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.640 0.000 10.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.640 0.000 10.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.640 0.000 10.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.640 0.000 10.792 0.152 ;
    END
  END O1[44]

  PIN I1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.424 0.000 9.576 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.424 0.000 9.576 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.424 0.000 9.576 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.424 0.000 9.576 0.152 ;
    END
  END I1[44]

  PIN I1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.120 0.000 9.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.120 0.000 9.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.120 0.000 9.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.120 0.000 9.272 0.152 ;
    END
  END I1[45]

  PIN I1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.816 0.000 8.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.816 0.000 8.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.816 0.000 8.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.816 0.000 8.968 0.152 ;
    END
  END I1[46]

  PIN I1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.512 0.000 8.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.512 0.000 8.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.512 0.000 8.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.512 0.000 8.664 0.152 ;
    END
  END I1[47]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.944 34.048 68.096 34.200 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.944 34.048 68.096 34.200 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.944 34.048 68.096 34.200 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.944 34.048 68.096 34.200 ;
    END
  END A1[0]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.944 30.400 68.096 30.552 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.944 30.400 68.096 30.552 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.944 30.400 68.096 30.552 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.944 30.400 68.096 30.552 ;
    END
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.944 26.752 68.096 26.904 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.944 26.752 68.096 26.904 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.944 26.752 68.096 26.904 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.944 26.752 68.096 26.904 ;
    END
  END A1[2]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.944 23.104 68.096 23.256 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.944 23.104 68.096 23.256 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.944 23.104 68.096 23.256 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.944 23.104 68.096 23.256 ;
    END
  END A1[3]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.944 19.456 68.096 19.608 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.944 19.456 68.096 19.608 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.944 19.456 68.096 19.608 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.944 19.456 68.096 19.608 ;
    END
  END A1[4]

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.944 15.808 68.096 15.960 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.944 15.808 68.096 15.960 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.944 15.808 68.096 15.960 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.944 15.808 68.096 15.960 ;
    END
  END A1[5]

  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.944 12.160 68.096 12.312 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.944 12.160 68.096 12.312 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.944 12.160 68.096 12.312 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.944 12.160 68.096 12.312 ;
    END
  END A1[6]

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.944 9.728 68.096 9.880 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.944 9.728 68.096 9.880 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.944 9.728 68.096 9.880 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.944 9.728 68.096 9.880 ;
    END
  END WEB1

  PIN WBM1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.944 8.512 68.096 8.664 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.944 8.512 68.096 8.664 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.944 8.512 68.096 8.664 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.944 8.512 68.096 8.664 ;
    END
  END WBM1[0]

  PIN WBM1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.944 7.296 68.096 7.448 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.944 7.296 68.096 7.448 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.944 7.296 68.096 7.448 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.944 7.296 68.096 7.448 ;
    END
  END WBM1[1]

  PIN WBM1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.944 6.080 68.096 6.232 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.944 6.080 68.096 6.232 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.944 6.080 68.096 6.232 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.944 6.080 68.096 6.232 ;
    END
  END WBM1[2]

  PIN WBM1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.944 4.864 68.096 5.016 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.944 4.864 68.096 5.016 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.944 4.864 68.096 5.016 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.944 4.864 68.096 5.016 ;
    END
  END WBM1[3]

  PIN WBM1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.944 3.648 68.096 3.800 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.944 3.648 68.096 3.800 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.944 3.648 68.096 3.800 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.944 3.648 68.096 3.800 ;
    END
  END WBM1[4]

  PIN WBM1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.944 2.432 68.096 2.584 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.944 2.432 68.096 2.584 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.944 2.432 68.096 2.584 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.944 2.432 68.096 2.584 ;
    END
  END WBM1[5]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 5.195 36.912 7.195 38.912 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.195 36.912 7.195 38.912 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.195 36.912 7.195 38.912 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M2 ;
        RECT 7.915 36.912 9.915 38.912 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.915 36.912 9.915 38.912 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.915 36.912 9.915 38.912 ;
    END
  END VSS

  OBS
    LAYER M2 ;
      RECT 62.320 0.000 68.096 0.304 ;
      RECT 61.104 0.000 61.864 0.304 ;
      RECT 59.888 0.000 60.648 0.304 ;
      RECT 58.672 0.000 59.432 0.304 ;
      RECT 56.544 0.000 57.304 0.304 ;
      RECT 54.416 0.000 55.176 0.304 ;
      RECT 52.288 0.000 53.048 0.304 ;
      RECT 50.160 0.000 50.920 0.304 ;
      RECT 48.032 0.000 48.792 0.304 ;
      RECT 45.904 0.000 46.664 0.304 ;
      RECT 43.776 0.000 44.536 0.304 ;
      RECT 41.648 0.000 42.408 0.304 ;
      RECT 39.520 0.000 40.280 0.304 ;
      RECT 37.392 0.000 38.152 0.304 ;
      RECT 35.264 0.000 36.024 0.304 ;
      RECT 33.136 0.000 33.896 0.304 ;
      RECT 31.008 0.000 31.768 0.304 ;
      RECT 28.880 0.000 29.640 0.304 ;
      RECT 26.752 0.000 27.512 0.304 ;
      RECT 24.624 0.000 25.384 0.304 ;
      RECT 22.496 0.000 23.256 0.304 ;
      RECT 20.368 0.000 21.128 0.304 ;
      RECT 18.240 0.000 19.000 0.304 ;
      RECT 16.112 0.000 16.872 0.304 ;
      RECT 13.984 0.000 14.744 0.304 ;
      RECT 11.856 0.000 12.616 0.304 ;
      RECT 9.728 0.000 10.488 0.304 ;
      RECT 0.000 0.000 8.360 0.304 ;
      RECT 67.792 34.352 68.096 36.760 ;
      RECT 67.792 30.704 68.096 33.896 ;
      RECT 67.792 27.056 68.096 30.248 ;
      RECT 67.792 23.408 68.096 26.600 ;
      RECT 67.792 19.760 68.096 22.952 ;
      RECT 67.792 16.112 68.096 19.304 ;
      RECT 67.792 12.464 68.096 15.656 ;
      RECT 67.792 10.032 68.096 12.008 ;
      RECT 67.792 8.816 68.096 9.576 ;
      RECT 67.792 7.600 68.096 8.360 ;
      RECT 67.792 6.384 68.096 7.144 ;
      RECT 67.792 5.168 68.096 5.928 ;
      RECT 67.792 3.952 68.096 4.712 ;
      RECT 67.792 2.736 68.096 3.496 ;
      RECT 67.792 0.304 68.096 2.280 ;
      RECT 0.000 36.760 5.043 38.912 ;
      RECT 7.355 36.760 7.763 38.912 ;
      RECT 10.067 36.760 68.096 38.912 ;
      RECT 0.000 0.304 67.792 36.760 ;
    LAYER M3 ;
      RECT 62.320 0.000 68.096 0.304 ;
      RECT 61.104 0.000 61.864 0.304 ;
      RECT 59.888 0.000 60.648 0.304 ;
      RECT 58.672 0.000 59.432 0.304 ;
      RECT 56.544 0.000 57.304 0.304 ;
      RECT 54.416 0.000 55.176 0.304 ;
      RECT 52.288 0.000 53.048 0.304 ;
      RECT 50.160 0.000 50.920 0.304 ;
      RECT 48.032 0.000 48.792 0.304 ;
      RECT 45.904 0.000 46.664 0.304 ;
      RECT 43.776 0.000 44.536 0.304 ;
      RECT 41.648 0.000 42.408 0.304 ;
      RECT 39.520 0.000 40.280 0.304 ;
      RECT 37.392 0.000 38.152 0.304 ;
      RECT 35.264 0.000 36.024 0.304 ;
      RECT 33.136 0.000 33.896 0.304 ;
      RECT 31.008 0.000 31.768 0.304 ;
      RECT 28.880 0.000 29.640 0.304 ;
      RECT 26.752 0.000 27.512 0.304 ;
      RECT 24.624 0.000 25.384 0.304 ;
      RECT 22.496 0.000 23.256 0.304 ;
      RECT 20.368 0.000 21.128 0.304 ;
      RECT 18.240 0.000 19.000 0.304 ;
      RECT 16.112 0.000 16.872 0.304 ;
      RECT 13.984 0.000 14.744 0.304 ;
      RECT 11.856 0.000 12.616 0.304 ;
      RECT 9.728 0.000 10.488 0.304 ;
      RECT 0.000 0.000 8.360 0.304 ;
      RECT 67.792 34.352 68.096 36.760 ;
      RECT 67.792 30.704 68.096 33.896 ;
      RECT 67.792 27.056 68.096 30.248 ;
      RECT 67.792 23.408 68.096 26.600 ;
      RECT 67.792 19.760 68.096 22.952 ;
      RECT 67.792 16.112 68.096 19.304 ;
      RECT 67.792 12.464 68.096 15.656 ;
      RECT 67.792 10.032 68.096 12.008 ;
      RECT 67.792 8.816 68.096 9.576 ;
      RECT 67.792 7.600 68.096 8.360 ;
      RECT 67.792 6.384 68.096 7.144 ;
      RECT 67.792 5.168 68.096 5.928 ;
      RECT 67.792 3.952 68.096 4.712 ;
      RECT 67.792 2.736 68.096 3.496 ;
      RECT 67.792 0.304 68.096 2.280 ;
      RECT 0.000 36.760 5.043 38.912 ;
      RECT 7.355 36.760 7.763 38.912 ;
      RECT 10.067 36.760 68.096 38.912 ;
      RECT 0.000 0.304 67.792 36.760 ;
    LAYER M4 ;
      RECT 62.320 0.000 68.096 0.304 ;
      RECT 61.104 0.000 61.864 0.304 ;
      RECT 59.888 0.000 60.648 0.304 ;
      RECT 58.672 0.000 59.432 0.304 ;
      RECT 56.544 0.000 57.304 0.304 ;
      RECT 54.416 0.000 55.176 0.304 ;
      RECT 52.288 0.000 53.048 0.304 ;
      RECT 50.160 0.000 50.920 0.304 ;
      RECT 48.032 0.000 48.792 0.304 ;
      RECT 45.904 0.000 46.664 0.304 ;
      RECT 43.776 0.000 44.536 0.304 ;
      RECT 41.648 0.000 42.408 0.304 ;
      RECT 39.520 0.000 40.280 0.304 ;
      RECT 37.392 0.000 38.152 0.304 ;
      RECT 35.264 0.000 36.024 0.304 ;
      RECT 33.136 0.000 33.896 0.304 ;
      RECT 31.008 0.000 31.768 0.304 ;
      RECT 28.880 0.000 29.640 0.304 ;
      RECT 26.752 0.000 27.512 0.304 ;
      RECT 24.624 0.000 25.384 0.304 ;
      RECT 22.496 0.000 23.256 0.304 ;
      RECT 20.368 0.000 21.128 0.304 ;
      RECT 18.240 0.000 19.000 0.304 ;
      RECT 16.112 0.000 16.872 0.304 ;
      RECT 13.984 0.000 14.744 0.304 ;
      RECT 11.856 0.000 12.616 0.304 ;
      RECT 9.728 0.000 10.488 0.304 ;
      RECT 0.000 0.000 8.360 0.304 ;
      RECT 67.792 34.352 68.096 36.760 ;
      RECT 67.792 30.704 68.096 33.896 ;
      RECT 67.792 27.056 68.096 30.248 ;
      RECT 67.792 23.408 68.096 26.600 ;
      RECT 67.792 19.760 68.096 22.952 ;
      RECT 67.792 16.112 68.096 19.304 ;
      RECT 67.792 12.464 68.096 15.656 ;
      RECT 67.792 10.032 68.096 12.008 ;
      RECT 67.792 8.816 68.096 9.576 ;
      RECT 67.792 7.600 68.096 8.360 ;
      RECT 67.792 6.384 68.096 7.144 ;
      RECT 67.792 5.168 68.096 5.928 ;
      RECT 67.792 3.952 68.096 4.712 ;
      RECT 67.792 2.736 68.096 3.496 ;
      RECT 67.792 0.304 68.096 2.280 ;
      RECT 0.000 36.760 5.043 38.912 ;
      RECT 7.355 36.760 7.763 38.912 ;
      RECT 10.067 36.760 68.096 38.912 ;
      RECT 0.000 0.304 67.792 36.760 ;
    LAYER M5 ;
      RECT 62.320 0.000 68.096 0.304 ;
      RECT 61.104 0.000 61.864 0.304 ;
      RECT 59.888 0.000 60.648 0.304 ;
      RECT 58.672 0.000 59.432 0.304 ;
      RECT 56.544 0.000 57.304 0.304 ;
      RECT 54.416 0.000 55.176 0.304 ;
      RECT 52.288 0.000 53.048 0.304 ;
      RECT 50.160 0.000 50.920 0.304 ;
      RECT 48.032 0.000 48.792 0.304 ;
      RECT 45.904 0.000 46.664 0.304 ;
      RECT 43.776 0.000 44.536 0.304 ;
      RECT 41.648 0.000 42.408 0.304 ;
      RECT 39.520 0.000 40.280 0.304 ;
      RECT 37.392 0.000 38.152 0.304 ;
      RECT 35.264 0.000 36.024 0.304 ;
      RECT 33.136 0.000 33.896 0.304 ;
      RECT 31.008 0.000 31.768 0.304 ;
      RECT 28.880 0.000 29.640 0.304 ;
      RECT 26.752 0.000 27.512 0.304 ;
      RECT 24.624 0.000 25.384 0.304 ;
      RECT 22.496 0.000 23.256 0.304 ;
      RECT 20.368 0.000 21.128 0.304 ;
      RECT 18.240 0.000 19.000 0.304 ;
      RECT 16.112 0.000 16.872 0.304 ;
      RECT 13.984 0.000 14.744 0.304 ;
      RECT 11.856 0.000 12.616 0.304 ;
      RECT 9.728 0.000 10.488 0.304 ;
      RECT 0.000 0.000 8.360 0.304 ;
      RECT 67.792 34.352 68.096 36.760 ;
      RECT 67.792 30.704 68.096 33.896 ;
      RECT 67.792 27.056 68.096 30.248 ;
      RECT 67.792 23.408 68.096 26.600 ;
      RECT 67.792 19.760 68.096 22.952 ;
      RECT 67.792 16.112 68.096 19.304 ;
      RECT 67.792 12.464 68.096 15.656 ;
      RECT 67.792 10.032 68.096 12.008 ;
      RECT 67.792 8.816 68.096 9.576 ;
      RECT 67.792 7.600 68.096 8.360 ;
      RECT 67.792 6.384 68.096 7.144 ;
      RECT 67.792 5.168 68.096 5.928 ;
      RECT 67.792 3.952 68.096 4.712 ;
      RECT 67.792 2.736 68.096 3.496 ;
      RECT 67.792 0.304 68.096 2.280 ;
      RECT 0.000 36.760 5.043 38.912 ;
      RECT 7.355 36.760 7.763 38.912 ;
      RECT 10.067 36.760 68.096 38.912 ;
      RECT 0.000 0.304 67.792 36.760 ;
  END

END sram6t128x48

END LIBRARY
