VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram8t32x144
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 120.256 BY 113.088 ;
  SYMMETRY X Y R90 ;

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.480 0.000 112.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 112.480 0.000 112.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.480 0.000 112.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.480 0.000 112.632 0.152 ;
    END
  END CE1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.176 0.000 112.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 112.176 0.000 112.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.176 0.000 112.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.176 0.000 112.328 0.152 ;
    END
  END CSB1

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.872 0.000 112.024 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 111.872 0.000 112.024 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 111.872 0.000 112.024 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.872 0.000 112.024 0.152 ;
    END
  END OEB1

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.568 0.000 111.720 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 111.568 0.000 111.720 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 111.568 0.000 111.720 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.568 0.000 111.720 0.152 ;
    END
  END O1[3]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.264 0.000 111.416 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 111.264 0.000 111.416 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 111.264 0.000 111.416 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.264 0.000 111.416 0.152 ;
    END
  END O1[2]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.960 0.000 111.112 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.960 0.000 111.112 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.960 0.000 111.112 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.960 0.000 111.112 0.152 ;
    END
  END O1[1]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.656 0.000 110.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.656 0.000 110.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.656 0.000 110.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.656 0.000 110.808 0.152 ;
    END
  END O1[0]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.352 0.000 110.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.352 0.000 110.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.352 0.000 110.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.352 0.000 110.504 0.152 ;
    END
  END O1[7]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
  END O1[6]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.744 0.000 109.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.744 0.000 109.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.744 0.000 109.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.744 0.000 109.896 0.152 ;
    END
  END O1[5]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.440 0.000 109.592 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.440 0.000 109.592 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.440 0.000 109.592 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.440 0.000 109.592 0.152 ;
    END
  END O1[4]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.136 0.000 109.288 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.136 0.000 109.288 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.136 0.000 109.288 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.136 0.000 109.288 0.152 ;
    END
  END O1[11]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.832 0.000 108.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.832 0.000 108.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.832 0.000 108.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.832 0.000 108.984 0.152 ;
    END
  END O1[10]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.528 0.000 108.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.528 0.000 108.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.528 0.000 108.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.528 0.000 108.680 0.152 ;
    END
  END O1[9]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.224 0.000 108.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.224 0.000 108.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.224 0.000 108.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.224 0.000 108.376 0.152 ;
    END
  END O1[8]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.920 0.000 108.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.920 0.000 108.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.920 0.000 108.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.920 0.000 108.072 0.152 ;
    END
  END O1[15]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.616 0.000 107.768 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.616 0.000 107.768 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.616 0.000 107.768 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.616 0.000 107.768 0.152 ;
    END
  END O1[14]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.312 0.000 107.464 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.312 0.000 107.464 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.312 0.000 107.464 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.312 0.000 107.464 0.152 ;
    END
  END O1[13]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.008 0.000 107.160 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.008 0.000 107.160 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.008 0.000 107.160 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.008 0.000 107.160 0.152 ;
    END
  END O1[12]

  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.704 0.000 106.856 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 106.704 0.000 106.856 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 106.704 0.000 106.856 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.704 0.000 106.856 0.152 ;
    END
  END O1[19]

  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.400 0.000 106.552 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 106.400 0.000 106.552 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 106.400 0.000 106.552 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.400 0.000 106.552 0.152 ;
    END
  END O1[18]

  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.096 0.000 106.248 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 106.096 0.000 106.248 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 106.096 0.000 106.248 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.096 0.000 106.248 0.152 ;
    END
  END O1[17]

  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.792 0.000 105.944 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.792 0.000 105.944 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.792 0.000 105.944 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.792 0.000 105.944 0.152 ;
    END
  END O1[16]

  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.488 0.000 105.640 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.488 0.000 105.640 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.488 0.000 105.640 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.488 0.000 105.640 0.152 ;
    END
  END O1[23]

  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.184 0.000 105.336 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.184 0.000 105.336 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.184 0.000 105.336 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.184 0.000 105.336 0.152 ;
    END
  END O1[22]

  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.880 0.000 105.032 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.880 0.000 105.032 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.880 0.000 105.032 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.880 0.000 105.032 0.152 ;
    END
  END O1[21]

  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.576 0.000 104.728 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.576 0.000 104.728 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.576 0.000 104.728 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.576 0.000 104.728 0.152 ;
    END
  END O1[20]

  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.272 0.000 104.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.272 0.000 104.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.272 0.000 104.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.272 0.000 104.424 0.152 ;
    END
  END O1[27]

  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.968 0.000 104.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.968 0.000 104.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.968 0.000 104.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.968 0.000 104.120 0.152 ;
    END
  END O1[26]

  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.664 0.000 103.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.664 0.000 103.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.664 0.000 103.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.664 0.000 103.816 0.152 ;
    END
  END O1[25]

  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.360 0.000 103.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.360 0.000 103.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.360 0.000 103.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.360 0.000 103.512 0.152 ;
    END
  END O1[24]

  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.056 0.000 103.208 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.056 0.000 103.208 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.056 0.000 103.208 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.056 0.000 103.208 0.152 ;
    END
  END O1[31]

  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.752 0.000 102.904 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.752 0.000 102.904 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.752 0.000 102.904 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.752 0.000 102.904 0.152 ;
    END
  END O1[30]

  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.448 0.000 102.600 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.448 0.000 102.600 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.448 0.000 102.600 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.448 0.000 102.600 0.152 ;
    END
  END O1[29]

  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.144 0.000 102.296 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.144 0.000 102.296 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.144 0.000 102.296 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.144 0.000 102.296 0.152 ;
    END
  END O1[28]

  PIN O1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.840 0.000 101.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.840 0.000 101.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.840 0.000 101.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.840 0.000 101.992 0.152 ;
    END
  END O1[35]

  PIN O1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.536 0.000 101.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.536 0.000 101.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.536 0.000 101.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.536 0.000 101.688 0.152 ;
    END
  END O1[34]

  PIN O1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.232 0.000 101.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.232 0.000 101.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.232 0.000 101.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.232 0.000 101.384 0.152 ;
    END
  END O1[33]

  PIN O1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.928 0.000 101.080 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.928 0.000 101.080 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.928 0.000 101.080 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.928 0.000 101.080 0.152 ;
    END
  END O1[32]

  PIN O1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.624 0.000 100.776 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.624 0.000 100.776 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.624 0.000 100.776 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.624 0.000 100.776 0.152 ;
    END
  END O1[39]

  PIN O1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.320 0.000 100.472 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.320 0.000 100.472 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.320 0.000 100.472 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.320 0.000 100.472 0.152 ;
    END
  END O1[38]

  PIN O1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.016 0.000 100.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.016 0.000 100.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.016 0.000 100.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.016 0.000 100.168 0.152 ;
    END
  END O1[37]

  PIN O1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.712 0.000 99.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.712 0.000 99.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.712 0.000 99.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.712 0.000 99.864 0.152 ;
    END
  END O1[36]

  PIN O1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.408 0.000 99.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.408 0.000 99.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.408 0.000 99.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.408 0.000 99.560 0.152 ;
    END
  END O1[43]

  PIN O1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.104 0.000 99.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.104 0.000 99.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.104 0.000 99.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.104 0.000 99.256 0.152 ;
    END
  END O1[42]

  PIN O1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.800 0.000 98.952 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.800 0.000 98.952 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.800 0.000 98.952 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.800 0.000 98.952 0.152 ;
    END
  END O1[41]

  PIN O1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.496 0.000 98.648 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.496 0.000 98.648 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.496 0.000 98.648 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.496 0.000 98.648 0.152 ;
    END
  END O1[40]

  PIN O1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.192 0.000 98.344 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.192 0.000 98.344 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.192 0.000 98.344 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.192 0.000 98.344 0.152 ;
    END
  END O1[47]

  PIN O1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.888 0.000 98.040 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.888 0.000 98.040 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.888 0.000 98.040 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.888 0.000 98.040 0.152 ;
    END
  END O1[46]

  PIN O1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.584 0.000 97.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.584 0.000 97.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.584 0.000 97.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.584 0.000 97.736 0.152 ;
    END
  END O1[45]

  PIN O1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.280 0.000 97.432 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.280 0.000 97.432 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.280 0.000 97.432 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.280 0.000 97.432 0.152 ;
    END
  END O1[44]

  PIN O1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.976 0.000 97.128 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.976 0.000 97.128 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.976 0.000 97.128 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.976 0.000 97.128 0.152 ;
    END
  END O1[51]

  PIN O1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.672 0.000 96.824 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.672 0.000 96.824 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.672 0.000 96.824 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.672 0.000 96.824 0.152 ;
    END
  END O1[50]

  PIN O1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.368 0.000 96.520 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.368 0.000 96.520 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.368 0.000 96.520 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.368 0.000 96.520 0.152 ;
    END
  END O1[49]

  PIN O1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.064 0.000 96.216 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.064 0.000 96.216 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.064 0.000 96.216 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.064 0.000 96.216 0.152 ;
    END
  END O1[48]

  PIN O1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.760 0.000 95.912 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.760 0.000 95.912 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.760 0.000 95.912 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.760 0.000 95.912 0.152 ;
    END
  END O1[55]

  PIN O1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.456 0.000 95.608 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.456 0.000 95.608 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.456 0.000 95.608 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.456 0.000 95.608 0.152 ;
    END
  END O1[54]

  PIN O1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.152 0.000 95.304 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.152 0.000 95.304 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.152 0.000 95.304 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.152 0.000 95.304 0.152 ;
    END
  END O1[53]

  PIN O1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.848 0.000 95.000 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.848 0.000 95.000 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.848 0.000 95.000 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.848 0.000 95.000 0.152 ;
    END
  END O1[52]

  PIN O1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.544 0.000 94.696 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.544 0.000 94.696 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.544 0.000 94.696 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.544 0.000 94.696 0.152 ;
    END
  END O1[59]

  PIN O1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.240 0.000 94.392 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.240 0.000 94.392 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.240 0.000 94.392 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.240 0.000 94.392 0.152 ;
    END
  END O1[58]

  PIN O1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.936 0.000 94.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.936 0.000 94.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.936 0.000 94.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.936 0.000 94.088 0.152 ;
    END
  END O1[57]

  PIN O1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.632 0.000 93.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.632 0.000 93.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.632 0.000 93.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.632 0.000 93.784 0.152 ;
    END
  END O1[56]

  PIN O1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.328 0.000 93.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.328 0.000 93.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.328 0.000 93.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.328 0.000 93.480 0.152 ;
    END
  END O1[63]

  PIN O1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
  END O1[62]

  PIN O1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.720 0.000 92.872 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.720 0.000 92.872 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.720 0.000 92.872 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.720 0.000 92.872 0.152 ;
    END
  END O1[61]

  PIN O1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.416 0.000 92.568 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.416 0.000 92.568 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.416 0.000 92.568 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.416 0.000 92.568 0.152 ;
    END
  END O1[60]

  PIN O1[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.112 0.000 92.264 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.112 0.000 92.264 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.112 0.000 92.264 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.112 0.000 92.264 0.152 ;
    END
  END O1[67]

  PIN O1[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.808 0.000 91.960 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 91.808 0.000 91.960 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 91.808 0.000 91.960 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.808 0.000 91.960 0.152 ;
    END
  END O1[66]

  PIN O1[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.504 0.000 91.656 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 91.504 0.000 91.656 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 91.504 0.000 91.656 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.504 0.000 91.656 0.152 ;
    END
  END O1[65]

  PIN O1[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.200 0.000 91.352 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 91.200 0.000 91.352 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 91.200 0.000 91.352 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.200 0.000 91.352 0.152 ;
    END
  END O1[64]

  PIN O1[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.896 0.000 91.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.896 0.000 91.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.896 0.000 91.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.896 0.000 91.048 0.152 ;
    END
  END O1[71]

  PIN O1[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.592 0.000 90.744 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.592 0.000 90.744 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.592 0.000 90.744 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.592 0.000 90.744 0.152 ;
    END
  END O1[70]

  PIN O1[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.288 0.000 90.440 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.288 0.000 90.440 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.288 0.000 90.440 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.288 0.000 90.440 0.152 ;
    END
  END O1[69]

  PIN O1[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.984 0.000 90.136 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.984 0.000 90.136 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.984 0.000 90.136 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.984 0.000 90.136 0.152 ;
    END
  END O1[68]

  PIN O1[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.680 0.000 89.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.680 0.000 89.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.680 0.000 89.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.680 0.000 89.832 0.152 ;
    END
  END O1[75]

  PIN O1[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.376 0.000 89.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.376 0.000 89.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.376 0.000 89.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.376 0.000 89.528 0.152 ;
    END
  END O1[74]

  PIN O1[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.072 0.000 89.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.072 0.000 89.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.072 0.000 89.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.072 0.000 89.224 0.152 ;
    END
  END O1[73]

  PIN O1[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
  END O1[72]

  PIN O1[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
  END O1[79]

  PIN O1[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
  END O1[78]

  PIN O1[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
  END O1[77]

  PIN O1[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.552 0.000 87.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.552 0.000 87.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.552 0.000 87.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.552 0.000 87.704 0.152 ;
    END
  END O1[76]

  PIN O1[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.248 0.000 87.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.248 0.000 87.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.248 0.000 87.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.248 0.000 87.400 0.152 ;
    END
  END O1[83]

  PIN O1[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.944 0.000 87.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.944 0.000 87.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.944 0.000 87.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.944 0.000 87.096 0.152 ;
    END
  END O1[82]

  PIN O1[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.640 0.000 86.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.640 0.000 86.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.640 0.000 86.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.640 0.000 86.792 0.152 ;
    END
  END O1[81]

  PIN O1[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.336 0.000 86.488 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.336 0.000 86.488 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.336 0.000 86.488 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.336 0.000 86.488 0.152 ;
    END
  END O1[80]

  PIN O1[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.032 0.000 86.184 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.032 0.000 86.184 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.032 0.000 86.184 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.032 0.000 86.184 0.152 ;
    END
  END O1[87]

  PIN O1[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.728 0.000 85.880 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.728 0.000 85.880 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.728 0.000 85.880 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.728 0.000 85.880 0.152 ;
    END
  END O1[86]

  PIN O1[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.424 0.000 85.576 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.424 0.000 85.576 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.424 0.000 85.576 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.424 0.000 85.576 0.152 ;
    END
  END O1[85]

  PIN O1[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.120 0.000 85.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.120 0.000 85.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.120 0.000 85.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.120 0.000 85.272 0.152 ;
    END
  END O1[84]

  PIN O1[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.816 0.000 84.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.816 0.000 84.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.816 0.000 84.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.816 0.000 84.968 0.152 ;
    END
  END O1[91]

  PIN O1[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.512 0.000 84.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.512 0.000 84.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.512 0.000 84.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.512 0.000 84.664 0.152 ;
    END
  END O1[90]

  PIN O1[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.208 0.000 84.360 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.208 0.000 84.360 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.208 0.000 84.360 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.208 0.000 84.360 0.152 ;
    END
  END O1[89]

  PIN O1[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.904 0.000 84.056 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.904 0.000 84.056 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.904 0.000 84.056 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.904 0.000 84.056 0.152 ;
    END
  END O1[88]

  PIN O1[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.600 0.000 83.752 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.600 0.000 83.752 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.600 0.000 83.752 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.600 0.000 83.752 0.152 ;
    END
  END O1[95]

  PIN O1[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.296 0.000 83.448 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.296 0.000 83.448 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.296 0.000 83.448 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.296 0.000 83.448 0.152 ;
    END
  END O1[94]

  PIN O1[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.992 0.000 83.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.992 0.000 83.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.992 0.000 83.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.992 0.000 83.144 0.152 ;
    END
  END O1[93]

  PIN O1[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.688 0.000 82.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.688 0.000 82.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.688 0.000 82.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.688 0.000 82.840 0.152 ;
    END
  END O1[92]

  PIN O1[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
  END O1[99]

  PIN O1[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.080 0.000 82.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.080 0.000 82.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.080 0.000 82.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.080 0.000 82.232 0.152 ;
    END
  END O1[98]

  PIN O1[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.776 0.000 81.928 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.776 0.000 81.928 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.776 0.000 81.928 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.776 0.000 81.928 0.152 ;
    END
  END O1[97]

  PIN O1[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.472 0.000 81.624 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.472 0.000 81.624 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.472 0.000 81.624 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.472 0.000 81.624 0.152 ;
    END
  END O1[96]

  PIN O1[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.168 0.000 81.320 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.168 0.000 81.320 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.168 0.000 81.320 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.168 0.000 81.320 0.152 ;
    END
  END O1[103]

  PIN O1[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.864 0.000 81.016 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.864 0.000 81.016 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.864 0.000 81.016 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.864 0.000 81.016 0.152 ;
    END
  END O1[102]

  PIN O1[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.560 0.000 80.712 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.560 0.000 80.712 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.560 0.000 80.712 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.560 0.000 80.712 0.152 ;
    END
  END O1[101]

  PIN O1[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.256 0.000 80.408 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.256 0.000 80.408 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.256 0.000 80.408 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.256 0.000 80.408 0.152 ;
    END
  END O1[100]

  PIN O1[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.952 0.000 80.104 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.952 0.000 80.104 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.952 0.000 80.104 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.952 0.000 80.104 0.152 ;
    END
  END O1[107]

  PIN O1[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.648 0.000 79.800 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.648 0.000 79.800 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.648 0.000 79.800 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.648 0.000 79.800 0.152 ;
    END
  END O1[106]

  PIN O1[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.344 0.000 79.496 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.344 0.000 79.496 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.344 0.000 79.496 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.344 0.000 79.496 0.152 ;
    END
  END O1[105]

  PIN O1[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.040 0.000 79.192 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.040 0.000 79.192 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.040 0.000 79.192 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.040 0.000 79.192 0.152 ;
    END
  END O1[104]

  PIN O1[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.736 0.000 78.888 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.736 0.000 78.888 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.736 0.000 78.888 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.736 0.000 78.888 0.152 ;
    END
  END O1[111]

  PIN O1[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.432 0.000 78.584 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.432 0.000 78.584 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.432 0.000 78.584 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.432 0.000 78.584 0.152 ;
    END
  END O1[110]

  PIN O1[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.128 0.000 78.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.128 0.000 78.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.128 0.000 78.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.128 0.000 78.280 0.152 ;
    END
  END O1[109]

  PIN O1[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.824 0.000 77.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.824 0.000 77.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.824 0.000 77.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.824 0.000 77.976 0.152 ;
    END
  END O1[108]

  PIN O1[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.520 0.000 77.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.520 0.000 77.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.520 0.000 77.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.520 0.000 77.672 0.152 ;
    END
  END O1[115]

  PIN O1[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.216 0.000 77.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.216 0.000 77.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.216 0.000 77.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.216 0.000 77.368 0.152 ;
    END
  END O1[114]

  PIN O1[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.912 0.000 77.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.912 0.000 77.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.912 0.000 77.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.912 0.000 77.064 0.152 ;
    END
  END O1[113]

  PIN O1[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.608 0.000 76.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.608 0.000 76.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.608 0.000 76.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.608 0.000 76.760 0.152 ;
    END
  END O1[112]

  PIN O1[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.304 0.000 76.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.304 0.000 76.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.304 0.000 76.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.304 0.000 76.456 0.152 ;
    END
  END O1[119]

  PIN O1[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.000 0.000 76.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.000 0.000 76.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.000 0.000 76.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.000 0.000 76.152 0.152 ;
    END
  END O1[118]

  PIN O1[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.696 0.000 75.848 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.696 0.000 75.848 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.696 0.000 75.848 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.696 0.000 75.848 0.152 ;
    END
  END O1[117]

  PIN O1[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.392 0.000 75.544 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.392 0.000 75.544 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.392 0.000 75.544 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.392 0.000 75.544 0.152 ;
    END
  END O1[116]

  PIN O1[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.088 0.000 75.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.088 0.000 75.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.088 0.000 75.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.088 0.000 75.240 0.152 ;
    END
  END O1[123]

  PIN O1[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.784 0.000 74.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.784 0.000 74.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.784 0.000 74.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.784 0.000 74.936 0.152 ;
    END
  END O1[122]

  PIN O1[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.480 0.000 74.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.480 0.000 74.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.480 0.000 74.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.480 0.000 74.632 0.152 ;
    END
  END O1[121]

  PIN O1[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.176 0.000 74.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.176 0.000 74.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.176 0.000 74.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.176 0.000 74.328 0.152 ;
    END
  END O1[120]

  PIN O1[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.872 0.000 74.024 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.872 0.000 74.024 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.872 0.000 74.024 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.872 0.000 74.024 0.152 ;
    END
  END O1[127]

  PIN O1[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.568 0.000 73.720 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.568 0.000 73.720 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.568 0.000 73.720 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.568 0.000 73.720 0.152 ;
    END
  END O1[126]

  PIN O1[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.264 0.000 73.416 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.264 0.000 73.416 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.264 0.000 73.416 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.264 0.000 73.416 0.152 ;
    END
  END O1[125]

  PIN O1[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.960 0.000 73.112 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.960 0.000 73.112 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.960 0.000 73.112 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.960 0.000 73.112 0.152 ;
    END
  END O1[124]

  PIN O1[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.656 0.000 72.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.656 0.000 72.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.656 0.000 72.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.656 0.000 72.808 0.152 ;
    END
  END O1[131]

  PIN O1[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.352 0.000 72.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.352 0.000 72.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.352 0.000 72.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.352 0.000 72.504 0.152 ;
    END
  END O1[130]

  PIN O1[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.048 0.000 72.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.048 0.000 72.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.048 0.000 72.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.048 0.000 72.200 0.152 ;
    END
  END O1[129]

  PIN O1[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
  END O1[128]

  PIN O1[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.440 0.000 71.592 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.440 0.000 71.592 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.440 0.000 71.592 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.440 0.000 71.592 0.152 ;
    END
  END O1[135]

  PIN O1[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.136 0.000 71.288 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.136 0.000 71.288 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.136 0.000 71.288 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.136 0.000 71.288 0.152 ;
    END
  END O1[134]

  PIN O1[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.832 0.000 70.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.832 0.000 70.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.832 0.000 70.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.832 0.000 70.984 0.152 ;
    END
  END O1[133]

  PIN O1[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.528 0.000 70.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.528 0.000 70.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.528 0.000 70.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.528 0.000 70.680 0.152 ;
    END
  END O1[132]

  PIN O1[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.224 0.000 70.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.224 0.000 70.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.224 0.000 70.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.224 0.000 70.376 0.152 ;
    END
  END O1[139]

  PIN O1[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.920 0.000 70.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.920 0.000 70.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.920 0.000 70.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.920 0.000 70.072 0.152 ;
    END
  END O1[138]

  PIN O1[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.616 0.000 69.768 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.616 0.000 69.768 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.616 0.000 69.768 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.616 0.000 69.768 0.152 ;
    END
  END O1[137]

  PIN O1[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.312 0.000 69.464 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.312 0.000 69.464 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.312 0.000 69.464 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.312 0.000 69.464 0.152 ;
    END
  END O1[136]

  PIN O1[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.008 0.000 69.160 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.008 0.000 69.160 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.008 0.000 69.160 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.008 0.000 69.160 0.152 ;
    END
  END O1[143]

  PIN O1[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.704 0.000 68.856 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.704 0.000 68.856 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.704 0.000 68.856 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.704 0.000 68.856 0.152 ;
    END
  END O1[142]

  PIN O1[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.400 0.000 68.552 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.400 0.000 68.552 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.400 0.000 68.552 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.400 0.000 68.552 0.152 ;
    END
  END O1[141]

  PIN O1[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.096 0.000 68.248 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.096 0.000 68.248 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.096 0.000 68.248 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.096 0.000 68.248 0.152 ;
    END
  END O1[140]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.104 98.952 120.256 99.104 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.104 98.952 120.256 99.104 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.104 98.952 120.256 99.104 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.104 98.952 120.256 99.104 ;
    END
  END A1[0]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.104 95.304 120.256 95.456 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.104 95.304 120.256 95.456 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.104 95.304 120.256 95.456 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.104 95.304 120.256 95.456 ;
    END
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.104 91.656 120.256 91.808 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.104 91.656 120.256 91.808 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.104 91.656 120.256 91.808 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.104 91.656 120.256 91.808 ;
    END
  END A1[2]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.104 88.008 120.256 88.160 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.104 88.008 120.256 88.160 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.104 88.008 120.256 88.160 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.104 88.008 120.256 88.160 ;
    END
  END A1[3]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.104 84.360 120.256 84.512 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.104 84.360 120.256 84.512 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.104 84.360 120.256 84.512 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.104 84.360 120.256 84.512 ;
    END
  END A1[4]

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 7.776 0.000 7.928 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.776 0.000 7.928 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 7.776 0.000 7.928 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.776 0.000 7.928 0.152 ;
    END
  END CE2

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.080 0.000 8.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.080 0.000 8.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.080 0.000 8.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.080 0.000 8.232 0.152 ;
    END
  END CSB2

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.384 0.000 8.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.384 0.000 8.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.384 0.000 8.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.384 0.000 8.536 0.152 ;
    END
  END I2[0]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.688 0.000 8.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.688 0.000 8.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.688 0.000 8.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.688 0.000 8.840 0.152 ;
    END
  END I2[1]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.992 0.000 9.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 8.992 0.000 9.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.992 0.000 9.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 8.992 0.000 9.144 0.152 ;
    END
  END I2[2]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.296 0.000 9.448 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.296 0.000 9.448 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.296 0.000 9.448 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.296 0.000 9.448 0.152 ;
    END
  END I2[3]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.600 0.000 9.752 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.600 0.000 9.752 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.600 0.000 9.752 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.600 0.000 9.752 0.152 ;
    END
  END I2[4]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.904 0.000 10.056 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.904 0.000 10.056 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.904 0.000 10.056 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.904 0.000 10.056 0.152 ;
    END
  END I2[5]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.208 0.000 10.360 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.208 0.000 10.360 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.208 0.000 10.360 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.208 0.000 10.360 0.152 ;
    END
  END I2[6]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.512 0.000 10.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.512 0.000 10.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.512 0.000 10.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.512 0.000 10.664 0.152 ;
    END
  END I2[7]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.816 0.000 10.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.816 0.000 10.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.816 0.000 10.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.816 0.000 10.968 0.152 ;
    END
  END I2[8]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.120 0.000 11.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.120 0.000 11.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.120 0.000 11.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.120 0.000 11.272 0.152 ;
    END
  END I2[9]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.424 0.000 11.576 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.424 0.000 11.576 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.424 0.000 11.576 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.424 0.000 11.576 0.152 ;
    END
  END I2[10]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.728 0.000 11.880 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.728 0.000 11.880 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.728 0.000 11.880 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.728 0.000 11.880 0.152 ;
    END
  END I2[11]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.032 0.000 12.184 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.032 0.000 12.184 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.032 0.000 12.184 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.032 0.000 12.184 0.152 ;
    END
  END I2[12]

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.336 0.000 12.488 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.336 0.000 12.488 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.336 0.000 12.488 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.336 0.000 12.488 0.152 ;
    END
  END I2[13]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.640 0.000 12.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.640 0.000 12.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.640 0.000 12.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.640 0.000 12.792 0.152 ;
    END
  END I2[14]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.944 0.000 13.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 12.944 0.000 13.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 12.944 0.000 13.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 12.944 0.000 13.096 0.152 ;
    END
  END I2[15]

  PIN I2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.248 0.000 13.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.248 0.000 13.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.248 0.000 13.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.248 0.000 13.400 0.152 ;
    END
  END I2[16]

  PIN I2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.552 0.000 13.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.552 0.000 13.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.552 0.000 13.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.552 0.000 13.704 0.152 ;
    END
  END I2[17]

  PIN I2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.856 0.000 14.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.856 0.000 14.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.856 0.000 14.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.856 0.000 14.008 0.152 ;
    END
  END I2[18]

  PIN I2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.160 0.000 14.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 14.160 0.000 14.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 14.160 0.000 14.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.160 0.000 14.312 0.152 ;
    END
  END I2[19]

  PIN I2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.464 0.000 14.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 14.464 0.000 14.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 14.464 0.000 14.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.464 0.000 14.616 0.152 ;
    END
  END I2[20]

  PIN I2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.768 0.000 14.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 14.768 0.000 14.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 14.768 0.000 14.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.768 0.000 14.920 0.152 ;
    END
  END I2[21]

  PIN I2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.072 0.000 15.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.072 0.000 15.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.072 0.000 15.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.072 0.000 15.224 0.152 ;
    END
  END I2[22]

  PIN I2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.376 0.000 15.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.376 0.000 15.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.376 0.000 15.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.376 0.000 15.528 0.152 ;
    END
  END I2[23]

  PIN I2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.680 0.000 15.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.680 0.000 15.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.680 0.000 15.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.680 0.000 15.832 0.152 ;
    END
  END I2[24]

  PIN I2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.984 0.000 16.136 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.984 0.000 16.136 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.984 0.000 16.136 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.984 0.000 16.136 0.152 ;
    END
  END I2[25]

  PIN I2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.288 0.000 16.440 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.288 0.000 16.440 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.288 0.000 16.440 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.288 0.000 16.440 0.152 ;
    END
  END I2[26]

  PIN I2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.592 0.000 16.744 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.592 0.000 16.744 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.592 0.000 16.744 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.592 0.000 16.744 0.152 ;
    END
  END I2[27]

  PIN I2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.896 0.000 17.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.896 0.000 17.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.896 0.000 17.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.896 0.000 17.048 0.152 ;
    END
  END I2[28]

  PIN I2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.200 0.000 17.352 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.200 0.000 17.352 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.200 0.000 17.352 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.200 0.000 17.352 0.152 ;
    END
  END I2[29]

  PIN I2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.504 0.000 17.656 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.504 0.000 17.656 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.504 0.000 17.656 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.504 0.000 17.656 0.152 ;
    END
  END I2[30]

  PIN I2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.808 0.000 17.960 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.808 0.000 17.960 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.808 0.000 17.960 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.808 0.000 17.960 0.152 ;
    END
  END I2[31]

  PIN I2[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.112 0.000 18.264 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.112 0.000 18.264 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.112 0.000 18.264 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.112 0.000 18.264 0.152 ;
    END
  END I2[32]

  PIN I2[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.416 0.000 18.568 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.416 0.000 18.568 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.416 0.000 18.568 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.416 0.000 18.568 0.152 ;
    END
  END I2[33]

  PIN I2[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.720 0.000 18.872 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 18.720 0.000 18.872 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 18.720 0.000 18.872 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 18.720 0.000 18.872 0.152 ;
    END
  END I2[34]

  PIN I2[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.024 0.000 19.176 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.024 0.000 19.176 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.024 0.000 19.176 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.024 0.000 19.176 0.152 ;
    END
  END I2[35]

  PIN I2[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.328 0.000 19.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.328 0.000 19.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.328 0.000 19.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.328 0.000 19.480 0.152 ;
    END
  END I2[36]

  PIN I2[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.632 0.000 19.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.632 0.000 19.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.632 0.000 19.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.632 0.000 19.784 0.152 ;
    END
  END I2[37]

  PIN I2[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.936 0.000 20.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.936 0.000 20.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.936 0.000 20.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.936 0.000 20.088 0.152 ;
    END
  END I2[38]

  PIN I2[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.240 0.000 20.392 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.240 0.000 20.392 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.240 0.000 20.392 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.240 0.000 20.392 0.152 ;
    END
  END I2[39]

  PIN I2[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.544 0.000 20.696 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.544 0.000 20.696 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.544 0.000 20.696 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.544 0.000 20.696 0.152 ;
    END
  END I2[40]

  PIN I2[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.848 0.000 21.000 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.848 0.000 21.000 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.848 0.000 21.000 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.848 0.000 21.000 0.152 ;
    END
  END I2[41]

  PIN I2[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.152 0.000 21.304 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.152 0.000 21.304 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.152 0.000 21.304 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.152 0.000 21.304 0.152 ;
    END
  END I2[42]

  PIN I2[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.456 0.000 21.608 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.456 0.000 21.608 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.456 0.000 21.608 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.456 0.000 21.608 0.152 ;
    END
  END I2[43]

  PIN I2[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.760 0.000 21.912 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.760 0.000 21.912 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.760 0.000 21.912 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.760 0.000 21.912 0.152 ;
    END
  END I2[44]

  PIN I2[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.064 0.000 22.216 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.064 0.000 22.216 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.064 0.000 22.216 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.064 0.000 22.216 0.152 ;
    END
  END I2[45]

  PIN I2[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.368 0.000 22.520 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.368 0.000 22.520 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.368 0.000 22.520 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.368 0.000 22.520 0.152 ;
    END
  END I2[46]

  PIN I2[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.672 0.000 22.824 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.672 0.000 22.824 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.672 0.000 22.824 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.672 0.000 22.824 0.152 ;
    END
  END I2[47]

  PIN I2[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.976 0.000 23.128 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.976 0.000 23.128 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.976 0.000 23.128 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.976 0.000 23.128 0.152 ;
    END
  END I2[48]

  PIN I2[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.280 0.000 23.432 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.280 0.000 23.432 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.280 0.000 23.432 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.280 0.000 23.432 0.152 ;
    END
  END I2[49]

  PIN I2[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.584 0.000 23.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.584 0.000 23.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.584 0.000 23.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.584 0.000 23.736 0.152 ;
    END
  END I2[50]

  PIN I2[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.888 0.000 24.040 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.888 0.000 24.040 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.888 0.000 24.040 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.888 0.000 24.040 0.152 ;
    END
  END I2[51]

  PIN I2[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.192 0.000 24.344 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.192 0.000 24.344 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.192 0.000 24.344 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.192 0.000 24.344 0.152 ;
    END
  END I2[52]

  PIN I2[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.496 0.000 24.648 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.496 0.000 24.648 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.496 0.000 24.648 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.496 0.000 24.648 0.152 ;
    END
  END I2[53]

  PIN I2[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.800 0.000 24.952 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.800 0.000 24.952 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.800 0.000 24.952 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.800 0.000 24.952 0.152 ;
    END
  END I2[54]

  PIN I2[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.104 0.000 25.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.104 0.000 25.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.104 0.000 25.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.104 0.000 25.256 0.152 ;
    END
  END I2[55]

  PIN I2[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.408 0.000 25.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.408 0.000 25.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.408 0.000 25.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.408 0.000 25.560 0.152 ;
    END
  END I2[56]

  PIN I2[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.712 0.000 25.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.712 0.000 25.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.712 0.000 25.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.712 0.000 25.864 0.152 ;
    END
  END I2[57]

  PIN I2[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.016 0.000 26.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.016 0.000 26.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.016 0.000 26.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.016 0.000 26.168 0.152 ;
    END
  END I2[58]

  PIN I2[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.320 0.000 26.472 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.320 0.000 26.472 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.320 0.000 26.472 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.320 0.000 26.472 0.152 ;
    END
  END I2[59]

  PIN I2[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.624 0.000 26.776 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.624 0.000 26.776 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.624 0.000 26.776 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.624 0.000 26.776 0.152 ;
    END
  END I2[60]

  PIN I2[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.928 0.000 27.080 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.928 0.000 27.080 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.928 0.000 27.080 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.928 0.000 27.080 0.152 ;
    END
  END I2[61]

  PIN I2[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.232 0.000 27.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.232 0.000 27.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.232 0.000 27.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.232 0.000 27.384 0.152 ;
    END
  END I2[62]

  PIN I2[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.536 0.000 27.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.536 0.000 27.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.536 0.000 27.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.536 0.000 27.688 0.152 ;
    END
  END I2[63]

  PIN I2[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.840 0.000 27.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.840 0.000 27.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.840 0.000 27.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.840 0.000 27.992 0.152 ;
    END
  END I2[64]

  PIN I2[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.144 0.000 28.296 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.144 0.000 28.296 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.144 0.000 28.296 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.144 0.000 28.296 0.152 ;
    END
  END I2[65]

  PIN I2[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.448 0.000 28.600 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.448 0.000 28.600 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.448 0.000 28.600 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.448 0.000 28.600 0.152 ;
    END
  END I2[66]

  PIN I2[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.752 0.000 28.904 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.752 0.000 28.904 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.752 0.000 28.904 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.752 0.000 28.904 0.152 ;
    END
  END I2[67]

  PIN I2[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.056 0.000 29.208 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.056 0.000 29.208 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.056 0.000 29.208 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.056 0.000 29.208 0.152 ;
    END
  END I2[68]

  PIN I2[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.360 0.000 29.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.360 0.000 29.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.360 0.000 29.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.360 0.000 29.512 0.152 ;
    END
  END I2[69]

  PIN I2[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.664 0.000 29.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.664 0.000 29.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.664 0.000 29.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.664 0.000 29.816 0.152 ;
    END
  END I2[70]

  PIN I2[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.968 0.000 30.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.968 0.000 30.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.968 0.000 30.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.968 0.000 30.120 0.152 ;
    END
  END I2[71]

  PIN I2[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.272 0.000 30.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.272 0.000 30.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.272 0.000 30.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.272 0.000 30.424 0.152 ;
    END
  END I2[72]

  PIN I2[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.576 0.000 30.728 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.576 0.000 30.728 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.576 0.000 30.728 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.576 0.000 30.728 0.152 ;
    END
  END I2[73]

  PIN I2[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.880 0.000 31.032 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.880 0.000 31.032 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.880 0.000 31.032 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.880 0.000 31.032 0.152 ;
    END
  END I2[74]

  PIN I2[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.184 0.000 31.336 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.184 0.000 31.336 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.184 0.000 31.336 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.184 0.000 31.336 0.152 ;
    END
  END I2[75]

  PIN I2[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.488 0.000 31.640 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.488 0.000 31.640 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.488 0.000 31.640 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.488 0.000 31.640 0.152 ;
    END
  END I2[76]

  PIN I2[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.792 0.000 31.944 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.792 0.000 31.944 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.792 0.000 31.944 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.792 0.000 31.944 0.152 ;
    END
  END I2[77]

  PIN I2[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.096 0.000 32.248 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.096 0.000 32.248 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.096 0.000 32.248 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.096 0.000 32.248 0.152 ;
    END
  END I2[78]

  PIN I2[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.400 0.000 32.552 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.400 0.000 32.552 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.400 0.000 32.552 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.400 0.000 32.552 0.152 ;
    END
  END I2[79]

  PIN I2[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.704 0.000 32.856 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.704 0.000 32.856 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.704 0.000 32.856 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.704 0.000 32.856 0.152 ;
    END
  END I2[80]

  PIN I2[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.008 0.000 33.160 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.008 0.000 33.160 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.008 0.000 33.160 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.008 0.000 33.160 0.152 ;
    END
  END I2[81]

  PIN I2[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.312 0.000 33.464 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.312 0.000 33.464 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.312 0.000 33.464 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.312 0.000 33.464 0.152 ;
    END
  END I2[82]

  PIN I2[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.616 0.000 33.768 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.616 0.000 33.768 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.616 0.000 33.768 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.616 0.000 33.768 0.152 ;
    END
  END I2[83]

  PIN I2[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.920 0.000 34.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.920 0.000 34.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.920 0.000 34.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.920 0.000 34.072 0.152 ;
    END
  END I2[84]

  PIN I2[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.224 0.000 34.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.224 0.000 34.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.224 0.000 34.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.224 0.000 34.376 0.152 ;
    END
  END I2[85]

  PIN I2[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.528 0.000 34.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.528 0.000 34.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.528 0.000 34.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.528 0.000 34.680 0.152 ;
    END
  END I2[86]

  PIN I2[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.832 0.000 34.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.832 0.000 34.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.832 0.000 34.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.832 0.000 34.984 0.152 ;
    END
  END I2[87]

  PIN I2[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.136 0.000 35.288 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.136 0.000 35.288 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.136 0.000 35.288 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.136 0.000 35.288 0.152 ;
    END
  END I2[88]

  PIN I2[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.440 0.000 35.592 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.440 0.000 35.592 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.440 0.000 35.592 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.440 0.000 35.592 0.152 ;
    END
  END I2[89]

  PIN I2[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.744 0.000 35.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.744 0.000 35.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.744 0.000 35.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.744 0.000 35.896 0.152 ;
    END
  END I2[90]

  PIN I2[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.048 0.000 36.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.048 0.000 36.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.048 0.000 36.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.048 0.000 36.200 0.152 ;
    END
  END I2[91]

  PIN I2[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.352 0.000 36.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.352 0.000 36.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.352 0.000 36.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.352 0.000 36.504 0.152 ;
    END
  END I2[92]

  PIN I2[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.656 0.000 36.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.656 0.000 36.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.656 0.000 36.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.656 0.000 36.808 0.152 ;
    END
  END I2[93]

  PIN I2[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.960 0.000 37.112 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.960 0.000 37.112 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.960 0.000 37.112 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.960 0.000 37.112 0.152 ;
    END
  END I2[94]

  PIN I2[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.264 0.000 37.416 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.264 0.000 37.416 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.264 0.000 37.416 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.264 0.000 37.416 0.152 ;
    END
  END I2[95]

  PIN I2[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.568 0.000 37.720 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.568 0.000 37.720 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.568 0.000 37.720 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.568 0.000 37.720 0.152 ;
    END
  END I2[96]

  PIN I2[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.872 0.000 38.024 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.872 0.000 38.024 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.872 0.000 38.024 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.872 0.000 38.024 0.152 ;
    END
  END I2[97]

  PIN I2[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.176 0.000 38.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.176 0.000 38.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.176 0.000 38.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.176 0.000 38.328 0.152 ;
    END
  END I2[98]

  PIN I2[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.480 0.000 38.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.480 0.000 38.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.480 0.000 38.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.480 0.000 38.632 0.152 ;
    END
  END I2[99]

  PIN I2[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.784 0.000 38.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.784 0.000 38.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.784 0.000 38.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.784 0.000 38.936 0.152 ;
    END
  END I2[100]

  PIN I2[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.088 0.000 39.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.088 0.000 39.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.088 0.000 39.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.088 0.000 39.240 0.152 ;
    END
  END I2[101]

  PIN I2[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.392 0.000 39.544 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.392 0.000 39.544 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.392 0.000 39.544 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.392 0.000 39.544 0.152 ;
    END
  END I2[102]

  PIN I2[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.696 0.000 39.848 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.696 0.000 39.848 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.696 0.000 39.848 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.696 0.000 39.848 0.152 ;
    END
  END I2[103]

  PIN I2[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.000 0.000 40.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.000 0.000 40.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.000 0.000 40.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.000 0.000 40.152 0.152 ;
    END
  END I2[104]

  PIN I2[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.304 0.000 40.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.304 0.000 40.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.304 0.000 40.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.304 0.000 40.456 0.152 ;
    END
  END I2[105]

  PIN I2[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.608 0.000 40.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.608 0.000 40.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.608 0.000 40.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.608 0.000 40.760 0.152 ;
    END
  END I2[106]

  PIN I2[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.912 0.000 41.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.912 0.000 41.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.912 0.000 41.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.912 0.000 41.064 0.152 ;
    END
  END I2[107]

  PIN I2[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.216 0.000 41.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.216 0.000 41.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.216 0.000 41.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.216 0.000 41.368 0.152 ;
    END
  END I2[108]

  PIN I2[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.520 0.000 41.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.520 0.000 41.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.520 0.000 41.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.520 0.000 41.672 0.152 ;
    END
  END I2[109]

  PIN I2[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.824 0.000 41.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.824 0.000 41.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.824 0.000 41.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.824 0.000 41.976 0.152 ;
    END
  END I2[110]

  PIN I2[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.128 0.000 42.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.128 0.000 42.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.128 0.000 42.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.128 0.000 42.280 0.152 ;
    END
  END I2[111]

  PIN I2[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.432 0.000 42.584 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.432 0.000 42.584 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.432 0.000 42.584 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.432 0.000 42.584 0.152 ;
    END
  END I2[112]

  PIN I2[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.736 0.000 42.888 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.736 0.000 42.888 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.736 0.000 42.888 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.736 0.000 42.888 0.152 ;
    END
  END I2[113]

  PIN I2[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.040 0.000 43.192 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.040 0.000 43.192 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.040 0.000 43.192 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.040 0.000 43.192 0.152 ;
    END
  END I2[114]

  PIN I2[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.344 0.000 43.496 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.344 0.000 43.496 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.344 0.000 43.496 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.344 0.000 43.496 0.152 ;
    END
  END I2[115]

  PIN I2[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.648 0.000 43.800 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.648 0.000 43.800 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.648 0.000 43.800 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.648 0.000 43.800 0.152 ;
    END
  END I2[116]

  PIN I2[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.952 0.000 44.104 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.952 0.000 44.104 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.952 0.000 44.104 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.952 0.000 44.104 0.152 ;
    END
  END I2[117]

  PIN I2[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.256 0.000 44.408 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.256 0.000 44.408 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.256 0.000 44.408 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.256 0.000 44.408 0.152 ;
    END
  END I2[118]

  PIN I2[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.560 0.000 44.712 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.560 0.000 44.712 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.560 0.000 44.712 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.560 0.000 44.712 0.152 ;
    END
  END I2[119]

  PIN I2[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.864 0.000 45.016 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.864 0.000 45.016 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.864 0.000 45.016 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.864 0.000 45.016 0.152 ;
    END
  END I2[120]

  PIN I2[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.168 0.000 45.320 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.168 0.000 45.320 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.168 0.000 45.320 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.168 0.000 45.320 0.152 ;
    END
  END I2[121]

  PIN I2[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.472 0.000 45.624 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.472 0.000 45.624 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.472 0.000 45.624 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.472 0.000 45.624 0.152 ;
    END
  END I2[122]

  PIN I2[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.776 0.000 45.928 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.776 0.000 45.928 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.776 0.000 45.928 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.776 0.000 45.928 0.152 ;
    END
  END I2[123]

  PIN I2[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.080 0.000 46.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.080 0.000 46.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.080 0.000 46.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.080 0.000 46.232 0.152 ;
    END
  END I2[124]

  PIN I2[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.384 0.000 46.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.384 0.000 46.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.384 0.000 46.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.384 0.000 46.536 0.152 ;
    END
  END I2[125]

  PIN I2[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.688 0.000 46.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.688 0.000 46.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.688 0.000 46.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.688 0.000 46.840 0.152 ;
    END
  END I2[126]

  PIN I2[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.992 0.000 47.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.992 0.000 47.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.992 0.000 47.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.992 0.000 47.144 0.152 ;
    END
  END I2[127]

  PIN I2[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.296 0.000 47.448 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.296 0.000 47.448 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.296 0.000 47.448 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.296 0.000 47.448 0.152 ;
    END
  END I2[128]

  PIN I2[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.600 0.000 47.752 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.600 0.000 47.752 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.600 0.000 47.752 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.600 0.000 47.752 0.152 ;
    END
  END I2[129]

  PIN I2[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.904 0.000 48.056 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.904 0.000 48.056 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.904 0.000 48.056 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.904 0.000 48.056 0.152 ;
    END
  END I2[130]

  PIN I2[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.208 0.000 48.360 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.208 0.000 48.360 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.208 0.000 48.360 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.208 0.000 48.360 0.152 ;
    END
  END I2[131]

  PIN I2[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.512 0.000 48.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.512 0.000 48.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.512 0.000 48.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.512 0.000 48.664 0.152 ;
    END
  END I2[132]

  PIN I2[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.816 0.000 48.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.816 0.000 48.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.816 0.000 48.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.816 0.000 48.968 0.152 ;
    END
  END I2[133]

  PIN I2[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.120 0.000 49.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.120 0.000 49.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.120 0.000 49.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.120 0.000 49.272 0.152 ;
    END
  END I2[134]

  PIN I2[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.424 0.000 49.576 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.424 0.000 49.576 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.424 0.000 49.576 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.424 0.000 49.576 0.152 ;
    END
  END I2[135]

  PIN I2[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.728 0.000 49.880 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.728 0.000 49.880 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.728 0.000 49.880 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.728 0.000 49.880 0.152 ;
    END
  END I2[136]

  PIN I2[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.032 0.000 50.184 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.032 0.000 50.184 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.032 0.000 50.184 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.032 0.000 50.184 0.152 ;
    END
  END I2[137]

  PIN I2[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.336 0.000 50.488 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.336 0.000 50.488 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.336 0.000 50.488 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.336 0.000 50.488 0.152 ;
    END
  END I2[138]

  PIN I2[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.640 0.000 50.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.640 0.000 50.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.640 0.000 50.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.640 0.000 50.792 0.152 ;
    END
  END I2[139]

  PIN I2[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.944 0.000 51.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.944 0.000 51.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.944 0.000 51.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.944 0.000 51.096 0.152 ;
    END
  END I2[140]

  PIN I2[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.248 0.000 51.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.248 0.000 51.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.248 0.000 51.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.248 0.000 51.400 0.152 ;
    END
  END I2[141]

  PIN I2[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.552 0.000 51.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.552 0.000 51.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.552 0.000 51.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.552 0.000 51.704 0.152 ;
    END
  END I2[142]

  PIN I2[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.856 0.000 52.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.856 0.000 52.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.856 0.000 52.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.856 0.000 52.008 0.152 ;
    END
  END I2[143]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 98.952 0.152 99.104 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 98.952 0.152 99.104 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 98.952 0.152 99.104 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 98.952 0.152 99.104 ;
    END
  END A2[0]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 95.304 0.152 95.456 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 95.304 0.152 95.456 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 95.304 0.152 95.456 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 95.304 0.152 95.456 ;
    END
  END A2[1]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 91.656 0.152 91.808 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 91.656 0.152 91.808 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 91.656 0.152 91.808 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 91.656 0.152 91.808 ;
    END
  END A2[2]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 88.008 0.152 88.160 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 88.008 0.152 88.160 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 88.008 0.152 88.160 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 88.008 0.152 88.160 ;
    END
  END A2[3]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 84.360 0.152 84.512 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 84.360 0.152 84.512 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 84.360 0.152 84.512 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 84.360 0.152 84.512 ;
    END
  END A2[4]

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 28.272 0.152 28.424 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 28.272 0.152 28.424 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 28.272 0.152 28.424 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 28.272 0.152 28.424 ;
    END
  END WEB2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 5.195 111.088 7.195 113.088 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.195 111.088 7.195 113.088 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.195 111.088 7.195 113.088 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M2 ;
        RECT 7.915 111.088 9.915 113.088 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.915 111.088 9.915 113.088 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.915 111.088 9.915 113.088 ;
    END
  END VSS

  OBS
    LAYER M2 ;
      RECT 112.784 0.000 120.256 0.304 ;
      RECT 112.480 0.000 112.328 0.304 ;
      RECT 112.176 0.000 112.024 0.304 ;
      RECT 111.872 0.000 111.720 0.304 ;
      RECT 110.656 0.000 110.504 0.304 ;
      RECT 109.440 0.000 109.288 0.304 ;
      RECT 108.224 0.000 108.072 0.304 ;
      RECT 107.008 0.000 106.856 0.304 ;
      RECT 105.792 0.000 105.640 0.304 ;
      RECT 104.576 0.000 104.424 0.304 ;
      RECT 103.360 0.000 103.208 0.304 ;
      RECT 102.144 0.000 101.992 0.304 ;
      RECT 100.928 0.000 100.776 0.304 ;
      RECT 99.712 0.000 99.560 0.304 ;
      RECT 98.496 0.000 98.344 0.304 ;
      RECT 97.280 0.000 97.128 0.304 ;
      RECT 96.064 0.000 95.912 0.304 ;
      RECT 94.848 0.000 94.696 0.304 ;
      RECT 93.632 0.000 93.480 0.304 ;
      RECT 92.416 0.000 92.264 0.304 ;
      RECT 91.200 0.000 91.048 0.304 ;
      RECT 89.984 0.000 89.832 0.304 ;
      RECT 88.768 0.000 88.616 0.304 ;
      RECT 87.552 0.000 87.400 0.304 ;
      RECT 86.336 0.000 86.184 0.304 ;
      RECT 85.120 0.000 84.968 0.304 ;
      RECT 83.904 0.000 83.752 0.304 ;
      RECT 82.688 0.000 82.536 0.304 ;
      RECT 81.472 0.000 81.320 0.304 ;
      RECT 80.256 0.000 80.104 0.304 ;
      RECT 79.040 0.000 78.888 0.304 ;
      RECT 77.824 0.000 77.672 0.304 ;
      RECT 76.608 0.000 76.456 0.304 ;
      RECT 75.392 0.000 75.240 0.304 ;
      RECT 74.176 0.000 74.024 0.304 ;
      RECT 72.960 0.000 72.808 0.304 ;
      RECT 71.744 0.000 71.592 0.304 ;
      RECT 70.528 0.000 70.376 0.304 ;
      RECT 69.312 0.000 69.160 0.304 ;
      RECT 119.952 99.256 120.256 110.936 ;
      RECT 119.952 95.608 120.256 98.800 ;
      RECT 119.952 91.960 120.256 95.152 ;
      RECT 119.952 88.312 120.256 91.504 ;
      RECT 119.952 84.664 120.256 87.856 ;
      RECT 119.952 28.576 120.256 84.208 ;
      RECT 119.952 0.304 120.256 28.120 ;
      RECT 0.000 0.000 7.624 0.304 ;
      RECT 8.080 0.000 7.928 0.304 ;
      RECT 8.384 0.000 8.232 0.304 ;
      RECT 9.600 0.000 9.448 0.304 ;
      RECT 10.816 0.000 10.664 0.304 ;
      RECT 12.032 0.000 11.880 0.304 ;
      RECT 13.248 0.000 13.096 0.304 ;
      RECT 14.464 0.000 14.312 0.304 ;
      RECT 15.680 0.000 15.528 0.304 ;
      RECT 16.896 0.000 16.744 0.304 ;
      RECT 18.112 0.000 17.960 0.304 ;
      RECT 19.328 0.000 19.176 0.304 ;
      RECT 20.544 0.000 20.392 0.304 ;
      RECT 21.760 0.000 21.608 0.304 ;
      RECT 22.976 0.000 22.824 0.304 ;
      RECT 24.192 0.000 24.040 0.304 ;
      RECT 25.408 0.000 25.256 0.304 ;
      RECT 26.624 0.000 26.472 0.304 ;
      RECT 27.840 0.000 27.688 0.304 ;
      RECT 29.056 0.000 28.904 0.304 ;
      RECT 30.272 0.000 30.120 0.304 ;
      RECT 31.488 0.000 31.336 0.304 ;
      RECT 32.704 0.000 32.552 0.304 ;
      RECT 33.920 0.000 33.768 0.304 ;
      RECT 35.136 0.000 34.984 0.304 ;
      RECT 36.352 0.000 36.200 0.304 ;
      RECT 37.568 0.000 37.416 0.304 ;
      RECT 38.784 0.000 38.632 0.304 ;
      RECT 40.000 0.000 39.848 0.304 ;
      RECT 41.216 0.000 41.064 0.304 ;
      RECT 42.432 0.000 42.280 0.304 ;
      RECT 43.648 0.000 43.496 0.304 ;
      RECT 44.864 0.000 44.712 0.304 ;
      RECT 46.080 0.000 45.928 0.304 ;
      RECT 47.296 0.000 47.144 0.304 ;
      RECT 48.512 0.000 48.360 0.304 ;
      RECT 49.728 0.000 49.576 0.304 ;
      RECT 50.944 0.000 50.792 0.304 ;
      RECT 52.160 0.000 67.944 0.304 ;
      RECT 0.000 99.256 0.304 110.936 ;
      RECT 0.000 95.608 0.304 98.800 ;
      RECT 0.000 91.960 0.304 95.152 ;
      RECT 0.000 88.312 0.304 91.504 ;
      RECT 0.000 84.664 0.304 87.856 ;
      RECT 0.000 28.576 0.304 84.208 ;
      RECT 0.000 0.304 0.304 28.120 ;
      RECT 0.000 110.936 5.043 113.088 ;
      RECT 7.355 110.936 7.763 113.088 ;
      RECT 10.067 110.936 120.256 113.088 ;
      RECT 0.304 0.304 119.952 110.936 ;
    LAYER M3 ;
      RECT 112.784 0.000 120.256 0.304 ;
      RECT 112.480 0.000 112.328 0.304 ;
      RECT 112.176 0.000 112.024 0.304 ;
      RECT 111.872 0.000 111.720 0.304 ;
      RECT 110.656 0.000 110.504 0.304 ;
      RECT 109.440 0.000 109.288 0.304 ;
      RECT 108.224 0.000 108.072 0.304 ;
      RECT 107.008 0.000 106.856 0.304 ;
      RECT 105.792 0.000 105.640 0.304 ;
      RECT 104.576 0.000 104.424 0.304 ;
      RECT 103.360 0.000 103.208 0.304 ;
      RECT 102.144 0.000 101.992 0.304 ;
      RECT 100.928 0.000 100.776 0.304 ;
      RECT 99.712 0.000 99.560 0.304 ;
      RECT 98.496 0.000 98.344 0.304 ;
      RECT 97.280 0.000 97.128 0.304 ;
      RECT 96.064 0.000 95.912 0.304 ;
      RECT 94.848 0.000 94.696 0.304 ;
      RECT 93.632 0.000 93.480 0.304 ;
      RECT 92.416 0.000 92.264 0.304 ;
      RECT 91.200 0.000 91.048 0.304 ;
      RECT 89.984 0.000 89.832 0.304 ;
      RECT 88.768 0.000 88.616 0.304 ;
      RECT 87.552 0.000 87.400 0.304 ;
      RECT 86.336 0.000 86.184 0.304 ;
      RECT 85.120 0.000 84.968 0.304 ;
      RECT 83.904 0.000 83.752 0.304 ;
      RECT 82.688 0.000 82.536 0.304 ;
      RECT 81.472 0.000 81.320 0.304 ;
      RECT 80.256 0.000 80.104 0.304 ;
      RECT 79.040 0.000 78.888 0.304 ;
      RECT 77.824 0.000 77.672 0.304 ;
      RECT 76.608 0.000 76.456 0.304 ;
      RECT 75.392 0.000 75.240 0.304 ;
      RECT 74.176 0.000 74.024 0.304 ;
      RECT 72.960 0.000 72.808 0.304 ;
      RECT 71.744 0.000 71.592 0.304 ;
      RECT 70.528 0.000 70.376 0.304 ;
      RECT 69.312 0.000 69.160 0.304 ;
      RECT 119.952 99.256 120.256 110.936 ;
      RECT 119.952 95.608 120.256 98.800 ;
      RECT 119.952 91.960 120.256 95.152 ;
      RECT 119.952 88.312 120.256 91.504 ;
      RECT 119.952 84.664 120.256 87.856 ;
      RECT 119.952 28.576 120.256 84.208 ;
      RECT 119.952 0.304 120.256 28.120 ;
      RECT 0.000 0.000 7.624 0.304 ;
      RECT 8.080 0.000 7.928 0.304 ;
      RECT 8.384 0.000 8.232 0.304 ;
      RECT 9.600 0.000 9.448 0.304 ;
      RECT 10.816 0.000 10.664 0.304 ;
      RECT 12.032 0.000 11.880 0.304 ;
      RECT 13.248 0.000 13.096 0.304 ;
      RECT 14.464 0.000 14.312 0.304 ;
      RECT 15.680 0.000 15.528 0.304 ;
      RECT 16.896 0.000 16.744 0.304 ;
      RECT 18.112 0.000 17.960 0.304 ;
      RECT 19.328 0.000 19.176 0.304 ;
      RECT 20.544 0.000 20.392 0.304 ;
      RECT 21.760 0.000 21.608 0.304 ;
      RECT 22.976 0.000 22.824 0.304 ;
      RECT 24.192 0.000 24.040 0.304 ;
      RECT 25.408 0.000 25.256 0.304 ;
      RECT 26.624 0.000 26.472 0.304 ;
      RECT 27.840 0.000 27.688 0.304 ;
      RECT 29.056 0.000 28.904 0.304 ;
      RECT 30.272 0.000 30.120 0.304 ;
      RECT 31.488 0.000 31.336 0.304 ;
      RECT 32.704 0.000 32.552 0.304 ;
      RECT 33.920 0.000 33.768 0.304 ;
      RECT 35.136 0.000 34.984 0.304 ;
      RECT 36.352 0.000 36.200 0.304 ;
      RECT 37.568 0.000 37.416 0.304 ;
      RECT 38.784 0.000 38.632 0.304 ;
      RECT 40.000 0.000 39.848 0.304 ;
      RECT 41.216 0.000 41.064 0.304 ;
      RECT 42.432 0.000 42.280 0.304 ;
      RECT 43.648 0.000 43.496 0.304 ;
      RECT 44.864 0.000 44.712 0.304 ;
      RECT 46.080 0.000 45.928 0.304 ;
      RECT 47.296 0.000 47.144 0.304 ;
      RECT 48.512 0.000 48.360 0.304 ;
      RECT 49.728 0.000 49.576 0.304 ;
      RECT 50.944 0.000 50.792 0.304 ;
      RECT 52.160 0.000 67.944 0.304 ;
      RECT 0.000 99.256 0.304 110.936 ;
      RECT 0.000 95.608 0.304 98.800 ;
      RECT 0.000 91.960 0.304 95.152 ;
      RECT 0.000 88.312 0.304 91.504 ;
      RECT 0.000 84.664 0.304 87.856 ;
      RECT 0.000 28.576 0.304 84.208 ;
      RECT 0.000 0.304 0.304 28.120 ;
      RECT 0.000 110.936 5.043 113.088 ;
      RECT 7.355 110.936 7.763 113.088 ;
      RECT 10.067 110.936 120.256 113.088 ;
      RECT 0.304 0.304 119.952 110.936 ;
    LAYER M4 ;
      RECT 112.784 0.000 120.256 0.304 ;
      RECT 112.480 0.000 112.328 0.304 ;
      RECT 112.176 0.000 112.024 0.304 ;
      RECT 111.872 0.000 111.720 0.304 ;
      RECT 110.656 0.000 110.504 0.304 ;
      RECT 109.440 0.000 109.288 0.304 ;
      RECT 108.224 0.000 108.072 0.304 ;
      RECT 107.008 0.000 106.856 0.304 ;
      RECT 105.792 0.000 105.640 0.304 ;
      RECT 104.576 0.000 104.424 0.304 ;
      RECT 103.360 0.000 103.208 0.304 ;
      RECT 102.144 0.000 101.992 0.304 ;
      RECT 100.928 0.000 100.776 0.304 ;
      RECT 99.712 0.000 99.560 0.304 ;
      RECT 98.496 0.000 98.344 0.304 ;
      RECT 97.280 0.000 97.128 0.304 ;
      RECT 96.064 0.000 95.912 0.304 ;
      RECT 94.848 0.000 94.696 0.304 ;
      RECT 93.632 0.000 93.480 0.304 ;
      RECT 92.416 0.000 92.264 0.304 ;
      RECT 91.200 0.000 91.048 0.304 ;
      RECT 89.984 0.000 89.832 0.304 ;
      RECT 88.768 0.000 88.616 0.304 ;
      RECT 87.552 0.000 87.400 0.304 ;
      RECT 86.336 0.000 86.184 0.304 ;
      RECT 85.120 0.000 84.968 0.304 ;
      RECT 83.904 0.000 83.752 0.304 ;
      RECT 82.688 0.000 82.536 0.304 ;
      RECT 81.472 0.000 81.320 0.304 ;
      RECT 80.256 0.000 80.104 0.304 ;
      RECT 79.040 0.000 78.888 0.304 ;
      RECT 77.824 0.000 77.672 0.304 ;
      RECT 76.608 0.000 76.456 0.304 ;
      RECT 75.392 0.000 75.240 0.304 ;
      RECT 74.176 0.000 74.024 0.304 ;
      RECT 72.960 0.000 72.808 0.304 ;
      RECT 71.744 0.000 71.592 0.304 ;
      RECT 70.528 0.000 70.376 0.304 ;
      RECT 69.312 0.000 69.160 0.304 ;
      RECT 119.952 99.256 120.256 110.936 ;
      RECT 119.952 95.608 120.256 98.800 ;
      RECT 119.952 91.960 120.256 95.152 ;
      RECT 119.952 88.312 120.256 91.504 ;
      RECT 119.952 84.664 120.256 87.856 ;
      RECT 119.952 28.576 120.256 84.208 ;
      RECT 119.952 0.304 120.256 28.120 ;
      RECT 0.000 0.000 7.624 0.304 ;
      RECT 8.080 0.000 7.928 0.304 ;
      RECT 8.384 0.000 8.232 0.304 ;
      RECT 9.600 0.000 9.448 0.304 ;
      RECT 10.816 0.000 10.664 0.304 ;
      RECT 12.032 0.000 11.880 0.304 ;
      RECT 13.248 0.000 13.096 0.304 ;
      RECT 14.464 0.000 14.312 0.304 ;
      RECT 15.680 0.000 15.528 0.304 ;
      RECT 16.896 0.000 16.744 0.304 ;
      RECT 18.112 0.000 17.960 0.304 ;
      RECT 19.328 0.000 19.176 0.304 ;
      RECT 20.544 0.000 20.392 0.304 ;
      RECT 21.760 0.000 21.608 0.304 ;
      RECT 22.976 0.000 22.824 0.304 ;
      RECT 24.192 0.000 24.040 0.304 ;
      RECT 25.408 0.000 25.256 0.304 ;
      RECT 26.624 0.000 26.472 0.304 ;
      RECT 27.840 0.000 27.688 0.304 ;
      RECT 29.056 0.000 28.904 0.304 ;
      RECT 30.272 0.000 30.120 0.304 ;
      RECT 31.488 0.000 31.336 0.304 ;
      RECT 32.704 0.000 32.552 0.304 ;
      RECT 33.920 0.000 33.768 0.304 ;
      RECT 35.136 0.000 34.984 0.304 ;
      RECT 36.352 0.000 36.200 0.304 ;
      RECT 37.568 0.000 37.416 0.304 ;
      RECT 38.784 0.000 38.632 0.304 ;
      RECT 40.000 0.000 39.848 0.304 ;
      RECT 41.216 0.000 41.064 0.304 ;
      RECT 42.432 0.000 42.280 0.304 ;
      RECT 43.648 0.000 43.496 0.304 ;
      RECT 44.864 0.000 44.712 0.304 ;
      RECT 46.080 0.000 45.928 0.304 ;
      RECT 47.296 0.000 47.144 0.304 ;
      RECT 48.512 0.000 48.360 0.304 ;
      RECT 49.728 0.000 49.576 0.304 ;
      RECT 50.944 0.000 50.792 0.304 ;
      RECT 52.160 0.000 67.944 0.304 ;
      RECT 0.000 99.256 0.304 110.936 ;
      RECT 0.000 95.608 0.304 98.800 ;
      RECT 0.000 91.960 0.304 95.152 ;
      RECT 0.000 88.312 0.304 91.504 ;
      RECT 0.000 84.664 0.304 87.856 ;
      RECT 0.000 28.576 0.304 84.208 ;
      RECT 0.000 0.304 0.304 28.120 ;
      RECT 0.000 110.936 5.043 113.088 ;
      RECT 7.355 110.936 7.763 113.088 ;
      RECT 10.067 110.936 120.256 113.088 ;
      RECT 0.304 0.304 119.952 110.936 ;
    LAYER M5 ;
      RECT 112.784 0.000 120.256 0.304 ;
      RECT 112.480 0.000 112.328 0.304 ;
      RECT 112.176 0.000 112.024 0.304 ;
      RECT 111.872 0.000 111.720 0.304 ;
      RECT 110.656 0.000 110.504 0.304 ;
      RECT 109.440 0.000 109.288 0.304 ;
      RECT 108.224 0.000 108.072 0.304 ;
      RECT 107.008 0.000 106.856 0.304 ;
      RECT 105.792 0.000 105.640 0.304 ;
      RECT 104.576 0.000 104.424 0.304 ;
      RECT 103.360 0.000 103.208 0.304 ;
      RECT 102.144 0.000 101.992 0.304 ;
      RECT 100.928 0.000 100.776 0.304 ;
      RECT 99.712 0.000 99.560 0.304 ;
      RECT 98.496 0.000 98.344 0.304 ;
      RECT 97.280 0.000 97.128 0.304 ;
      RECT 96.064 0.000 95.912 0.304 ;
      RECT 94.848 0.000 94.696 0.304 ;
      RECT 93.632 0.000 93.480 0.304 ;
      RECT 92.416 0.000 92.264 0.304 ;
      RECT 91.200 0.000 91.048 0.304 ;
      RECT 89.984 0.000 89.832 0.304 ;
      RECT 88.768 0.000 88.616 0.304 ;
      RECT 87.552 0.000 87.400 0.304 ;
      RECT 86.336 0.000 86.184 0.304 ;
      RECT 85.120 0.000 84.968 0.304 ;
      RECT 83.904 0.000 83.752 0.304 ;
      RECT 82.688 0.000 82.536 0.304 ;
      RECT 81.472 0.000 81.320 0.304 ;
      RECT 80.256 0.000 80.104 0.304 ;
      RECT 79.040 0.000 78.888 0.304 ;
      RECT 77.824 0.000 77.672 0.304 ;
      RECT 76.608 0.000 76.456 0.304 ;
      RECT 75.392 0.000 75.240 0.304 ;
      RECT 74.176 0.000 74.024 0.304 ;
      RECT 72.960 0.000 72.808 0.304 ;
      RECT 71.744 0.000 71.592 0.304 ;
      RECT 70.528 0.000 70.376 0.304 ;
      RECT 69.312 0.000 69.160 0.304 ;
      RECT 119.952 99.256 120.256 110.936 ;
      RECT 119.952 95.608 120.256 98.800 ;
      RECT 119.952 91.960 120.256 95.152 ;
      RECT 119.952 88.312 120.256 91.504 ;
      RECT 119.952 84.664 120.256 87.856 ;
      RECT 119.952 28.576 120.256 84.208 ;
      RECT 119.952 0.304 120.256 28.120 ;
      RECT 0.000 0.000 7.624 0.304 ;
      RECT 8.080 0.000 7.928 0.304 ;
      RECT 8.384 0.000 8.232 0.304 ;
      RECT 9.600 0.000 9.448 0.304 ;
      RECT 10.816 0.000 10.664 0.304 ;
      RECT 12.032 0.000 11.880 0.304 ;
      RECT 13.248 0.000 13.096 0.304 ;
      RECT 14.464 0.000 14.312 0.304 ;
      RECT 15.680 0.000 15.528 0.304 ;
      RECT 16.896 0.000 16.744 0.304 ;
      RECT 18.112 0.000 17.960 0.304 ;
      RECT 19.328 0.000 19.176 0.304 ;
      RECT 20.544 0.000 20.392 0.304 ;
      RECT 21.760 0.000 21.608 0.304 ;
      RECT 22.976 0.000 22.824 0.304 ;
      RECT 24.192 0.000 24.040 0.304 ;
      RECT 25.408 0.000 25.256 0.304 ;
      RECT 26.624 0.000 26.472 0.304 ;
      RECT 27.840 0.000 27.688 0.304 ;
      RECT 29.056 0.000 28.904 0.304 ;
      RECT 30.272 0.000 30.120 0.304 ;
      RECT 31.488 0.000 31.336 0.304 ;
      RECT 32.704 0.000 32.552 0.304 ;
      RECT 33.920 0.000 33.768 0.304 ;
      RECT 35.136 0.000 34.984 0.304 ;
      RECT 36.352 0.000 36.200 0.304 ;
      RECT 37.568 0.000 37.416 0.304 ;
      RECT 38.784 0.000 38.632 0.304 ;
      RECT 40.000 0.000 39.848 0.304 ;
      RECT 41.216 0.000 41.064 0.304 ;
      RECT 42.432 0.000 42.280 0.304 ;
      RECT 43.648 0.000 43.496 0.304 ;
      RECT 44.864 0.000 44.712 0.304 ;
      RECT 46.080 0.000 45.928 0.304 ;
      RECT 47.296 0.000 47.144 0.304 ;
      RECT 48.512 0.000 48.360 0.304 ;
      RECT 49.728 0.000 49.576 0.304 ;
      RECT 50.944 0.000 50.792 0.304 ;
      RECT 52.160 0.000 67.944 0.304 ;
      RECT 0.000 99.256 0.304 110.936 ;
      RECT 0.000 95.608 0.304 98.800 ;
      RECT 0.000 91.960 0.304 95.152 ;
      RECT 0.000 88.312 0.304 91.504 ;
      RECT 0.000 84.664 0.304 87.856 ;
      RECT 0.000 28.576 0.304 84.208 ;
      RECT 0.000 0.304 0.304 28.120 ;
      RECT 0.000 110.936 5.043 113.088 ;
      RECT 7.355 110.936 7.763 113.088 ;
      RECT 10.067 110.936 120.256 113.088 ;
      RECT 0.304 0.304 119.952 110.936 ;
  END

END sram8t32x144

END LIBRARY
