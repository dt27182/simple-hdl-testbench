VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram8t512x128
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 278.464 BY 136.192 ;
  SYMMETRY X Y R90 ;

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 268.128 0.000 268.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 268.128 0.000 268.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 268.128 0.000 268.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 268.128 0.000 268.280 0.152 ;
    END
  END CE1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 265.392 0.000 265.544 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 265.392 0.000 265.544 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 265.392 0.000 265.544 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 265.392 0.000 265.544 0.152 ;
    END
  END CSB1

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 262.656 0.000 262.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 262.656 0.000 262.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 262.656 0.000 262.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 262.656 0.000 262.808 0.152 ;
    END
  END OEB1

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 259.920 0.000 260.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 259.920 0.000 260.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 259.920 0.000 260.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 259.920 0.000 260.072 0.152 ;
    END
  END O1[3]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 259.616 0.000 259.768 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 259.616 0.000 259.768 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 259.616 0.000 259.768 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 259.616 0.000 259.768 0.152 ;
    END
  END O1[2]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 259.312 0.000 259.464 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 259.312 0.000 259.464 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 259.312 0.000 259.464 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 259.312 0.000 259.464 0.152 ;
    END
  END O1[1]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 259.008 0.000 259.160 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 259.008 0.000 259.160 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 259.008 0.000 259.160 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 259.008 0.000 259.160 0.152 ;
    END
  END O1[0]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 256.272 0.000 256.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 256.272 0.000 256.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 256.272 0.000 256.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 256.272 0.000 256.424 0.152 ;
    END
  END O1[7]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.968 0.000 256.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 255.968 0.000 256.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 255.968 0.000 256.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 255.968 0.000 256.120 0.152 ;
    END
  END O1[6]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.664 0.000 255.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 255.664 0.000 255.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 255.664 0.000 255.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 255.664 0.000 255.816 0.152 ;
    END
  END O1[5]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 255.360 0.000 255.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 255.360 0.000 255.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 255.360 0.000 255.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 255.360 0.000 255.512 0.152 ;
    END
  END O1[4]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 252.624 0.000 252.776 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 252.624 0.000 252.776 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 252.624 0.000 252.776 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 252.624 0.000 252.776 0.152 ;
    END
  END O1[11]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 252.320 0.000 252.472 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 252.320 0.000 252.472 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 252.320 0.000 252.472 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 252.320 0.000 252.472 0.152 ;
    END
  END O1[10]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 252.016 0.000 252.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 252.016 0.000 252.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 252.016 0.000 252.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 252.016 0.000 252.168 0.152 ;
    END
  END O1[9]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 251.712 0.000 251.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 251.712 0.000 251.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 251.712 0.000 251.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 251.712 0.000 251.864 0.152 ;
    END
  END O1[8]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 248.976 0.000 249.128 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 248.976 0.000 249.128 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 248.976 0.000 249.128 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 248.976 0.000 249.128 0.152 ;
    END
  END O1[15]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 248.672 0.000 248.824 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 248.672 0.000 248.824 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 248.672 0.000 248.824 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 248.672 0.000 248.824 0.152 ;
    END
  END O1[14]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 248.368 0.000 248.520 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 248.368 0.000 248.520 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 248.368 0.000 248.520 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 248.368 0.000 248.520 0.152 ;
    END
  END O1[13]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 248.064 0.000 248.216 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 248.064 0.000 248.216 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 248.064 0.000 248.216 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 248.064 0.000 248.216 0.152 ;
    END
  END O1[12]

  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 245.328 0.000 245.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 245.328 0.000 245.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 245.328 0.000 245.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 245.328 0.000 245.480 0.152 ;
    END
  END O1[19]

  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 245.024 0.000 245.176 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 245.024 0.000 245.176 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 245.024 0.000 245.176 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 245.024 0.000 245.176 0.152 ;
    END
  END O1[18]

  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 244.720 0.000 244.872 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 244.720 0.000 244.872 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 244.720 0.000 244.872 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 244.720 0.000 244.872 0.152 ;
    END
  END O1[17]

  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 244.416 0.000 244.568 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 244.416 0.000 244.568 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 244.416 0.000 244.568 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 244.416 0.000 244.568 0.152 ;
    END
  END O1[16]

  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 241.680 0.000 241.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 241.680 0.000 241.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 241.680 0.000 241.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 241.680 0.000 241.832 0.152 ;
    END
  END O1[23]

  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 241.376 0.000 241.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 241.376 0.000 241.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 241.376 0.000 241.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 241.376 0.000 241.528 0.152 ;
    END
  END O1[22]

  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 241.072 0.000 241.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 241.072 0.000 241.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 241.072 0.000 241.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 241.072 0.000 241.224 0.152 ;
    END
  END O1[21]

  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 240.768 0.000 240.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 240.768 0.000 240.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 240.768 0.000 240.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 240.768 0.000 240.920 0.152 ;
    END
  END O1[20]

  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 238.032 0.000 238.184 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 238.032 0.000 238.184 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 238.032 0.000 238.184 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 238.032 0.000 238.184 0.152 ;
    END
  END O1[27]

  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 237.728 0.000 237.880 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 237.728 0.000 237.880 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 237.728 0.000 237.880 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 237.728 0.000 237.880 0.152 ;
    END
  END O1[26]

  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 237.424 0.000 237.576 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 237.424 0.000 237.576 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 237.424 0.000 237.576 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 237.424 0.000 237.576 0.152 ;
    END
  END O1[25]

  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 237.120 0.000 237.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 237.120 0.000 237.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 237.120 0.000 237.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 237.120 0.000 237.272 0.152 ;
    END
  END O1[24]

  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 234.384 0.000 234.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 234.384 0.000 234.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 234.384 0.000 234.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 234.384 0.000 234.536 0.152 ;
    END
  END O1[31]

  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 234.080 0.000 234.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 234.080 0.000 234.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 234.080 0.000 234.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 234.080 0.000 234.232 0.152 ;
    END
  END O1[30]

  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 233.776 0.000 233.928 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 233.776 0.000 233.928 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 233.776 0.000 233.928 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 233.776 0.000 233.928 0.152 ;
    END
  END O1[29]

  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 233.472 0.000 233.624 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 233.472 0.000 233.624 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 233.472 0.000 233.624 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 233.472 0.000 233.624 0.152 ;
    END
  END O1[28]

  PIN O1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 230.736 0.000 230.888 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 230.736 0.000 230.888 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 230.736 0.000 230.888 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 230.736 0.000 230.888 0.152 ;
    END
  END O1[35]

  PIN O1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 230.432 0.000 230.584 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 230.432 0.000 230.584 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 230.432 0.000 230.584 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 230.432 0.000 230.584 0.152 ;
    END
  END O1[34]

  PIN O1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 230.128 0.000 230.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 230.128 0.000 230.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 230.128 0.000 230.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 230.128 0.000 230.280 0.152 ;
    END
  END O1[33]

  PIN O1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 229.824 0.000 229.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 229.824 0.000 229.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 229.824 0.000 229.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 229.824 0.000 229.976 0.152 ;
    END
  END O1[32]

  PIN O1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 227.088 0.000 227.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 227.088 0.000 227.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 227.088 0.000 227.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 227.088 0.000 227.240 0.152 ;
    END
  END O1[39]

  PIN O1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.784 0.000 226.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 226.784 0.000 226.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 226.784 0.000 226.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 226.784 0.000 226.936 0.152 ;
    END
  END O1[38]

  PIN O1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.480 0.000 226.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 226.480 0.000 226.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 226.480 0.000 226.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 226.480 0.000 226.632 0.152 ;
    END
  END O1[37]

  PIN O1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 226.176 0.000 226.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 226.176 0.000 226.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 226.176 0.000 226.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 226.176 0.000 226.328 0.152 ;
    END
  END O1[36]

  PIN O1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 223.440 0.000 223.592 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 223.440 0.000 223.592 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 223.440 0.000 223.592 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 223.440 0.000 223.592 0.152 ;
    END
  END O1[43]

  PIN O1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 223.136 0.000 223.288 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 223.136 0.000 223.288 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 223.136 0.000 223.288 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 223.136 0.000 223.288 0.152 ;
    END
  END O1[42]

  PIN O1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.832 0.000 222.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 222.832 0.000 222.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 222.832 0.000 222.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 222.832 0.000 222.984 0.152 ;
    END
  END O1[41]

  PIN O1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 222.528 0.000 222.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 222.528 0.000 222.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 222.528 0.000 222.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 222.528 0.000 222.680 0.152 ;
    END
  END O1[40]

  PIN O1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.792 0.000 219.944 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 219.792 0.000 219.944 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 219.792 0.000 219.944 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 219.792 0.000 219.944 0.152 ;
    END
  END O1[47]

  PIN O1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.488 0.000 219.640 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 219.488 0.000 219.640 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 219.488 0.000 219.640 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 219.488 0.000 219.640 0.152 ;
    END
  END O1[46]

  PIN O1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 219.184 0.000 219.336 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 219.184 0.000 219.336 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 219.184 0.000 219.336 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 219.184 0.000 219.336 0.152 ;
    END
  END O1[45]

  PIN O1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 218.880 0.000 219.032 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 218.880 0.000 219.032 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 218.880 0.000 219.032 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 218.880 0.000 219.032 0.152 ;
    END
  END O1[44]

  PIN O1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.144 0.000 216.296 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 216.144 0.000 216.296 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 216.144 0.000 216.296 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 216.144 0.000 216.296 0.152 ;
    END
  END O1[51]

  PIN O1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.840 0.000 215.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 215.840 0.000 215.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 215.840 0.000 215.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 215.840 0.000 215.992 0.152 ;
    END
  END O1[50]

  PIN O1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.536 0.000 215.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 215.536 0.000 215.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 215.536 0.000 215.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 215.536 0.000 215.688 0.152 ;
    END
  END O1[49]

  PIN O1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.232 0.000 215.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 215.232 0.000 215.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 215.232 0.000 215.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 215.232 0.000 215.384 0.152 ;
    END
  END O1[48]

  PIN O1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 212.496 0.000 212.648 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 212.496 0.000 212.648 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 212.496 0.000 212.648 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 212.496 0.000 212.648 0.152 ;
    END
  END O1[55]

  PIN O1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 212.192 0.000 212.344 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 212.192 0.000 212.344 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 212.192 0.000 212.344 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 212.192 0.000 212.344 0.152 ;
    END
  END O1[54]

  PIN O1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.888 0.000 212.040 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 211.888 0.000 212.040 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 211.888 0.000 212.040 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 211.888 0.000 212.040 0.152 ;
    END
  END O1[53]

  PIN O1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.584 0.000 211.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 211.584 0.000 211.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 211.584 0.000 211.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 211.584 0.000 211.736 0.152 ;
    END
  END O1[52]

  PIN O1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 208.848 0.000 209.000 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 208.848 0.000 209.000 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 208.848 0.000 209.000 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 208.848 0.000 209.000 0.152 ;
    END
  END O1[59]

  PIN O1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 208.544 0.000 208.696 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 208.544 0.000 208.696 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 208.544 0.000 208.696 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 208.544 0.000 208.696 0.152 ;
    END
  END O1[58]

  PIN O1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 208.240 0.000 208.392 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 208.240 0.000 208.392 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 208.240 0.000 208.392 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 208.240 0.000 208.392 0.152 ;
    END
  END O1[57]

  PIN O1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.936 0.000 208.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 207.936 0.000 208.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 207.936 0.000 208.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 207.936 0.000 208.088 0.152 ;
    END
  END O1[56]

  PIN O1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.200 0.000 205.352 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.200 0.000 205.352 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.200 0.000 205.352 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.200 0.000 205.352 0.152 ;
    END
  END O1[63]

  PIN O1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.896 0.000 205.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 204.896 0.000 205.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 204.896 0.000 205.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 204.896 0.000 205.048 0.152 ;
    END
  END O1[62]

  PIN O1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.592 0.000 204.744 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 204.592 0.000 204.744 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 204.592 0.000 204.744 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 204.592 0.000 204.744 0.152 ;
    END
  END O1[61]

  PIN O1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 204.288 0.000 204.440 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 204.288 0.000 204.440 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 204.288 0.000 204.440 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 204.288 0.000 204.440 0.152 ;
    END
  END O1[60]

  PIN O1[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 201.552 0.000 201.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 201.552 0.000 201.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 201.552 0.000 201.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 201.552 0.000 201.704 0.152 ;
    END
  END O1[67]

  PIN O1[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 201.248 0.000 201.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 201.248 0.000 201.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 201.248 0.000 201.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 201.248 0.000 201.400 0.152 ;
    END
  END O1[66]

  PIN O1[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 200.944 0.000 201.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 200.944 0.000 201.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 200.944 0.000 201.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 200.944 0.000 201.096 0.152 ;
    END
  END O1[65]

  PIN O1[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 200.640 0.000 200.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 200.640 0.000 200.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 200.640 0.000 200.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 200.640 0.000 200.792 0.152 ;
    END
  END O1[64]

  PIN O1[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 197.904 0.000 198.056 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.904 0.000 198.056 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.904 0.000 198.056 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 197.904 0.000 198.056 0.152 ;
    END
  END O1[71]

  PIN O1[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 197.600 0.000 197.752 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.600 0.000 197.752 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.600 0.000 197.752 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 197.600 0.000 197.752 0.152 ;
    END
  END O1[70]

  PIN O1[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 197.296 0.000 197.448 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 197.296 0.000 197.448 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 197.296 0.000 197.448 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 197.296 0.000 197.448 0.152 ;
    END
  END O1[69]

  PIN O1[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 196.992 0.000 197.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 196.992 0.000 197.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 196.992 0.000 197.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 196.992 0.000 197.144 0.152 ;
    END
  END O1[68]

  PIN O1[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.256 0.000 194.408 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 194.256 0.000 194.408 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 194.256 0.000 194.408 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 194.256 0.000 194.408 0.152 ;
    END
  END O1[75]

  PIN O1[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 193.952 0.000 194.104 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 193.952 0.000 194.104 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 193.952 0.000 194.104 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 193.952 0.000 194.104 0.152 ;
    END
  END O1[74]

  PIN O1[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 193.648 0.000 193.800 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 193.648 0.000 193.800 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 193.648 0.000 193.800 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 193.648 0.000 193.800 0.152 ;
    END
  END O1[73]

  PIN O1[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 193.344 0.000 193.496 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 193.344 0.000 193.496 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 193.344 0.000 193.496 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 193.344 0.000 193.496 0.152 ;
    END
  END O1[72]

  PIN O1[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
  END O1[79]

  PIN O1[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.304 0.000 190.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 190.304 0.000 190.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 190.304 0.000 190.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.304 0.000 190.456 0.152 ;
    END
  END O1[78]

  PIN O1[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.000 0.000 190.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 190.000 0.000 190.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 190.000 0.000 190.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.000 0.000 190.152 0.152 ;
    END
  END O1[77]

  PIN O1[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 189.696 0.000 189.848 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 189.696 0.000 189.848 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 189.696 0.000 189.848 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 189.696 0.000 189.848 0.152 ;
    END
  END O1[76]

  PIN O1[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.960 0.000 187.112 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 186.960 0.000 187.112 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 186.960 0.000 187.112 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 186.960 0.000 187.112 0.152 ;
    END
  END O1[83]

  PIN O1[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.656 0.000 186.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 186.656 0.000 186.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 186.656 0.000 186.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 186.656 0.000 186.808 0.152 ;
    END
  END O1[82]

  PIN O1[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.352 0.000 186.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 186.352 0.000 186.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 186.352 0.000 186.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 186.352 0.000 186.504 0.152 ;
    END
  END O1[81]

  PIN O1[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.048 0.000 186.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 186.048 0.000 186.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 186.048 0.000 186.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 186.048 0.000 186.200 0.152 ;
    END
  END O1[80]

  PIN O1[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.312 0.000 183.464 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 183.312 0.000 183.464 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 183.312 0.000 183.464 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 183.312 0.000 183.464 0.152 ;
    END
  END O1[87]

  PIN O1[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.008 0.000 183.160 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 183.008 0.000 183.160 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 183.008 0.000 183.160 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 183.008 0.000 183.160 0.152 ;
    END
  END O1[86]

  PIN O1[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 182.704 0.000 182.856 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 182.704 0.000 182.856 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 182.704 0.000 182.856 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 182.704 0.000 182.856 0.152 ;
    END
  END O1[85]

  PIN O1[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 182.400 0.000 182.552 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 182.400 0.000 182.552 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 182.400 0.000 182.552 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 182.400 0.000 182.552 0.152 ;
    END
  END O1[84]

  PIN O1[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.664 0.000 179.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 179.664 0.000 179.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 179.664 0.000 179.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 179.664 0.000 179.816 0.152 ;
    END
  END O1[91]

  PIN O1[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.360 0.000 179.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 179.360 0.000 179.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 179.360 0.000 179.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 179.360 0.000 179.512 0.152 ;
    END
  END O1[90]

  PIN O1[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.056 0.000 179.208 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 179.056 0.000 179.208 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 179.056 0.000 179.208 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 179.056 0.000 179.208 0.152 ;
    END
  END O1[89]

  PIN O1[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.752 0.000 178.904 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 178.752 0.000 178.904 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 178.752 0.000 178.904 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 178.752 0.000 178.904 0.152 ;
    END
  END O1[88]

  PIN O1[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.016 0.000 176.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 176.016 0.000 176.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 176.016 0.000 176.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 176.016 0.000 176.168 0.152 ;
    END
  END O1[95]

  PIN O1[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.712 0.000 175.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 175.712 0.000 175.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 175.712 0.000 175.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.712 0.000 175.864 0.152 ;
    END
  END O1[94]

  PIN O1[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.408 0.000 175.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 175.408 0.000 175.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 175.408 0.000 175.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.408 0.000 175.560 0.152 ;
    END
  END O1[93]

  PIN O1[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.104 0.000 175.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 175.104 0.000 175.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 175.104 0.000 175.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.104 0.000 175.256 0.152 ;
    END
  END O1[92]

  PIN O1[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 172.368 0.000 172.520 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 172.368 0.000 172.520 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 172.368 0.000 172.520 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 172.368 0.000 172.520 0.152 ;
    END
  END O1[99]

  PIN O1[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 172.064 0.000 172.216 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 172.064 0.000 172.216 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 172.064 0.000 172.216 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 172.064 0.000 172.216 0.152 ;
    END
  END O1[98]

  PIN O1[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.760 0.000 171.912 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 171.760 0.000 171.912 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 171.760 0.000 171.912 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 171.760 0.000 171.912 0.152 ;
    END
  END O1[97]

  PIN O1[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.456 0.000 171.608 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 171.456 0.000 171.608 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 171.456 0.000 171.608 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 171.456 0.000 171.608 0.152 ;
    END
  END O1[96]

  PIN O1[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.720 0.000 168.872 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 168.720 0.000 168.872 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 168.720 0.000 168.872 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 168.720 0.000 168.872 0.152 ;
    END
  END O1[103]

  PIN O1[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.416 0.000 168.568 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 168.416 0.000 168.568 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 168.416 0.000 168.568 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 168.416 0.000 168.568 0.152 ;
    END
  END O1[102]

  PIN O1[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.112 0.000 168.264 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 168.112 0.000 168.264 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 168.112 0.000 168.264 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 168.112 0.000 168.264 0.152 ;
    END
  END O1[101]

  PIN O1[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.808 0.000 167.960 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 167.808 0.000 167.960 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 167.808 0.000 167.960 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 167.808 0.000 167.960 0.152 ;
    END
  END O1[100]

  PIN O1[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.072 0.000 165.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 165.072 0.000 165.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 165.072 0.000 165.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 165.072 0.000 165.224 0.152 ;
    END
  END O1[107]

  PIN O1[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.768 0.000 164.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 164.768 0.000 164.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 164.768 0.000 164.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 164.768 0.000 164.920 0.152 ;
    END
  END O1[106]

  PIN O1[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.464 0.000 164.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 164.464 0.000 164.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 164.464 0.000 164.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 164.464 0.000 164.616 0.152 ;
    END
  END O1[105]

  PIN O1[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.160 0.000 164.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 164.160 0.000 164.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 164.160 0.000 164.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 164.160 0.000 164.312 0.152 ;
    END
  END O1[104]

  PIN O1[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.424 0.000 161.576 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 161.424 0.000 161.576 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 161.424 0.000 161.576 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.424 0.000 161.576 0.152 ;
    END
  END O1[111]

  PIN O1[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.120 0.000 161.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 161.120 0.000 161.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 161.120 0.000 161.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.120 0.000 161.272 0.152 ;
    END
  END O1[110]

  PIN O1[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.816 0.000 160.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 160.816 0.000 160.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 160.816 0.000 160.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 160.816 0.000 160.968 0.152 ;
    END
  END O1[109]

  PIN O1[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.512 0.000 160.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 160.512 0.000 160.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 160.512 0.000 160.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 160.512 0.000 160.664 0.152 ;
    END
  END O1[108]

  PIN O1[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.776 0.000 157.928 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 157.776 0.000 157.928 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 157.776 0.000 157.928 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 157.776 0.000 157.928 0.152 ;
    END
  END O1[115]

  PIN O1[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.472 0.000 157.624 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 157.472 0.000 157.624 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 157.472 0.000 157.624 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 157.472 0.000 157.624 0.152 ;
    END
  END O1[114]

  PIN O1[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.168 0.000 157.320 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 157.168 0.000 157.320 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 157.168 0.000 157.320 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 157.168 0.000 157.320 0.152 ;
    END
  END O1[113]

  PIN O1[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.864 0.000 157.016 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 156.864 0.000 157.016 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 156.864 0.000 157.016 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 156.864 0.000 157.016 0.152 ;
    END
  END O1[112]

  PIN O1[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
  END O1[119]

  PIN O1[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
  END O1[118]

  PIN O1[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
  END O1[117]

  PIN O1[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
  END O1[116]

  PIN O1[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.480 0.000 150.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.480 0.000 150.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.480 0.000 150.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 150.480 0.000 150.632 0.152 ;
    END
  END O1[123]

  PIN O1[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.176 0.000 150.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.176 0.000 150.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.176 0.000 150.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 150.176 0.000 150.328 0.152 ;
    END
  END O1[122]

  PIN O1[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.872 0.000 150.024 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 149.872 0.000 150.024 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 149.872 0.000 150.024 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 149.872 0.000 150.024 0.152 ;
    END
  END O1[121]

  PIN O1[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.568 0.000 149.720 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 149.568 0.000 149.720 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 149.568 0.000 149.720 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 149.568 0.000 149.720 0.152 ;
    END
  END O1[120]

  PIN O1[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.832 0.000 146.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 146.832 0.000 146.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 146.832 0.000 146.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.832 0.000 146.984 0.152 ;
    END
  END O1[127]

  PIN O1[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.528 0.000 146.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 146.528 0.000 146.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 146.528 0.000 146.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.528 0.000 146.680 0.152 ;
    END
  END O1[126]

  PIN O1[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.224 0.000 146.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 146.224 0.000 146.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 146.224 0.000 146.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.224 0.000 146.376 0.152 ;
    END
  END O1[125]

  PIN O1[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.920 0.000 146.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 145.920 0.000 146.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 145.920 0.000 146.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.920 0.000 146.072 0.152 ;
    END
  END O1[124]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 119.168 278.464 119.320 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 119.168 278.464 119.320 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 119.168 278.464 119.320 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 119.168 278.464 119.320 ;
    END
  END A1[0]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 115.520 278.464 115.672 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 115.520 278.464 115.672 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 115.520 278.464 115.672 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 115.520 278.464 115.672 ;
    END
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 111.872 278.464 112.024 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 111.872 278.464 112.024 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 111.872 278.464 112.024 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 111.872 278.464 112.024 ;
    END
  END A1[2]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 108.224 278.464 108.376 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 108.224 278.464 108.376 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 108.224 278.464 108.376 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 108.224 278.464 108.376 ;
    END
  END A1[3]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 104.576 278.464 104.728 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 104.576 278.464 104.728 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 104.576 278.464 104.728 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 104.576 278.464 104.728 ;
    END
  END A1[4]

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 100.928 278.464 101.080 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 100.928 278.464 101.080 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 100.928 278.464 101.080 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 100.928 278.464 101.080 ;
    END
  END A1[5]

  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 97.280 278.464 97.432 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 97.280 278.464 97.432 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 97.280 278.464 97.432 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 97.280 278.464 97.432 ;
    END
  END A1[6]

  PIN A1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 93.632 278.464 93.784 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 93.632 278.464 93.784 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 93.632 278.464 93.784 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 93.632 278.464 93.784 ;
    END
  END A1[7]

  PIN A1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 278.312 89.984 278.464 90.136 ;
    END
    PORT
      LAYER M3 ;
        RECT 278.312 89.984 278.464 90.136 ;
    END
    PORT
      LAYER M4 ;
        RECT 278.312 89.984 278.464 90.136 ;
    END
    PORT
      LAYER M5 ;
        RECT 278.312 89.984 278.464 90.136 ;
    END
  END A1[8]

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.336 0.000 10.488 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.336 0.000 10.488 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.336 0.000 10.488 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.336 0.000 10.488 0.152 ;
    END
  END CE2

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.072 0.000 13.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.072 0.000 13.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.072 0.000 13.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.072 0.000 13.224 0.152 ;
    END
  END CSB2

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.808 0.000 15.960 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 15.808 0.000 15.960 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 15.808 0.000 15.960 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 15.808 0.000 15.960 0.152 ;
    END
  END I2[0]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.112 0.000 16.264 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.112 0.000 16.264 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.112 0.000 16.264 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.112 0.000 16.264 0.152 ;
    END
  END I2[1]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.416 0.000 16.568 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.416 0.000 16.568 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.416 0.000 16.568 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.416 0.000 16.568 0.152 ;
    END
  END I2[2]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.720 0.000 16.872 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.720 0.000 16.872 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.720 0.000 16.872 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.720 0.000 16.872 0.152 ;
    END
  END I2[3]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.456 0.000 19.608 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.456 0.000 19.608 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.456 0.000 19.608 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.456 0.000 19.608 0.152 ;
    END
  END I2[4]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.760 0.000 19.912 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 19.760 0.000 19.912 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 19.760 0.000 19.912 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 19.760 0.000 19.912 0.152 ;
    END
  END I2[5]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.064 0.000 20.216 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.064 0.000 20.216 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.064 0.000 20.216 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.064 0.000 20.216 0.152 ;
    END
  END I2[6]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.368 0.000 20.520 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.368 0.000 20.520 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.368 0.000 20.520 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.368 0.000 20.520 0.152 ;
    END
  END I2[7]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.104 0.000 23.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.104 0.000 23.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.104 0.000 23.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.104 0.000 23.256 0.152 ;
    END
  END I2[8]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.408 0.000 23.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.408 0.000 23.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.408 0.000 23.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.408 0.000 23.560 0.152 ;
    END
  END I2[9]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.712 0.000 23.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.712 0.000 23.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.712 0.000 23.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.712 0.000 23.864 0.152 ;
    END
  END I2[10]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.016 0.000 24.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.016 0.000 24.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.016 0.000 24.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.016 0.000 24.168 0.152 ;
    END
  END I2[11]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.752 0.000 26.904 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 26.752 0.000 26.904 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 26.752 0.000 26.904 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 26.752 0.000 26.904 0.152 ;
    END
  END I2[12]

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.056 0.000 27.208 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.056 0.000 27.208 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.056 0.000 27.208 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.056 0.000 27.208 0.152 ;
    END
  END I2[13]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.360 0.000 27.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.360 0.000 27.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.360 0.000 27.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.360 0.000 27.512 0.152 ;
    END
  END I2[14]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.664 0.000 27.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.664 0.000 27.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.664 0.000 27.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.664 0.000 27.816 0.152 ;
    END
  END I2[15]

  PIN I2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.400 0.000 30.552 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.400 0.000 30.552 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.400 0.000 30.552 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.400 0.000 30.552 0.152 ;
    END
  END I2[16]

  PIN I2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.704 0.000 30.856 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.704 0.000 30.856 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.704 0.000 30.856 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.704 0.000 30.856 0.152 ;
    END
  END I2[17]

  PIN I2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.008 0.000 31.160 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.008 0.000 31.160 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.008 0.000 31.160 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.008 0.000 31.160 0.152 ;
    END
  END I2[18]

  PIN I2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.312 0.000 31.464 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.312 0.000 31.464 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.312 0.000 31.464 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.312 0.000 31.464 0.152 ;
    END
  END I2[19]

  PIN I2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
  END I2[20]

  PIN I2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
  END I2[21]

  PIN I2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.656 0.000 34.808 0.152 ;
    END
  END I2[22]

  PIN I2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.960 0.000 35.112 0.152 ;
    END
  END I2[23]

  PIN I2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
  END I2[24]

  PIN I2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
  END I2[25]

  PIN I2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
  END I2[26]

  PIN I2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
  END I2[27]

  PIN I2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.344 0.000 41.496 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.344 0.000 41.496 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.344 0.000 41.496 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.344 0.000 41.496 0.152 ;
    END
  END I2[28]

  PIN I2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.648 0.000 41.800 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.648 0.000 41.800 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.648 0.000 41.800 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.648 0.000 41.800 0.152 ;
    END
  END I2[29]

  PIN I2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.952 0.000 42.104 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.952 0.000 42.104 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.952 0.000 42.104 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.952 0.000 42.104 0.152 ;
    END
  END I2[30]

  PIN I2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.256 0.000 42.408 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.256 0.000 42.408 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.256 0.000 42.408 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.256 0.000 42.408 0.152 ;
    END
  END I2[31]

  PIN I2[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.992 0.000 45.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.992 0.000 45.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.992 0.000 45.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.992 0.000 45.144 0.152 ;
    END
  END I2[32]

  PIN I2[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.296 0.000 45.448 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.296 0.000 45.448 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.296 0.000 45.448 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.296 0.000 45.448 0.152 ;
    END
  END I2[33]

  PIN I2[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.600 0.000 45.752 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.600 0.000 45.752 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.600 0.000 45.752 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.600 0.000 45.752 0.152 ;
    END
  END I2[34]

  PIN I2[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.904 0.000 46.056 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 45.904 0.000 46.056 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 45.904 0.000 46.056 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 45.904 0.000 46.056 0.152 ;
    END
  END I2[35]

  PIN I2[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.640 0.000 48.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.640 0.000 48.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.640 0.000 48.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.640 0.000 48.792 0.152 ;
    END
  END I2[36]

  PIN I2[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.944 0.000 49.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.944 0.000 49.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.944 0.000 49.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.944 0.000 49.096 0.152 ;
    END
  END I2[37]

  PIN I2[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
  END I2[38]

  PIN I2[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
  END I2[39]

  PIN I2[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.288 0.000 52.440 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.288 0.000 52.440 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.288 0.000 52.440 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.288 0.000 52.440 0.152 ;
    END
  END I2[40]

  PIN I2[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.592 0.000 52.744 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.592 0.000 52.744 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.592 0.000 52.744 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.592 0.000 52.744 0.152 ;
    END
  END I2[41]

  PIN I2[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.896 0.000 53.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.896 0.000 53.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.896 0.000 53.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.896 0.000 53.048 0.152 ;
    END
  END I2[42]

  PIN I2[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.200 0.000 53.352 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.200 0.000 53.352 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.200 0.000 53.352 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.200 0.000 53.352 0.152 ;
    END
  END I2[43]

  PIN I2[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.936 0.000 56.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.936 0.000 56.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.936 0.000 56.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.936 0.000 56.088 0.152 ;
    END
  END I2[44]

  PIN I2[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.240 0.000 56.392 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.240 0.000 56.392 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.240 0.000 56.392 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.240 0.000 56.392 0.152 ;
    END
  END I2[45]

  PIN I2[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.544 0.000 56.696 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.544 0.000 56.696 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.544 0.000 56.696 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.544 0.000 56.696 0.152 ;
    END
  END I2[46]

  PIN I2[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.848 0.000 57.000 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.848 0.000 57.000 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.848 0.000 57.000 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.848 0.000 57.000 0.152 ;
    END
  END I2[47]

  PIN I2[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.584 0.000 59.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.584 0.000 59.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.584 0.000 59.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.584 0.000 59.736 0.152 ;
    END
  END I2[48]

  PIN I2[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.888 0.000 60.040 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.888 0.000 60.040 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.888 0.000 60.040 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.888 0.000 60.040 0.152 ;
    END
  END I2[49]

  PIN I2[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.192 0.000 60.344 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.192 0.000 60.344 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.192 0.000 60.344 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.192 0.000 60.344 0.152 ;
    END
  END I2[50]

  PIN I2[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.496 0.000 60.648 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.496 0.000 60.648 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.496 0.000 60.648 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.496 0.000 60.648 0.152 ;
    END
  END I2[51]

  PIN I2[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.232 0.000 63.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.232 0.000 63.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.232 0.000 63.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.232 0.000 63.384 0.152 ;
    END
  END I2[52]

  PIN I2[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.536 0.000 63.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.536 0.000 63.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.536 0.000 63.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.536 0.000 63.688 0.152 ;
    END
  END I2[53]

  PIN I2[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.840 0.000 63.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.840 0.000 63.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.840 0.000 63.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.840 0.000 63.992 0.152 ;
    END
  END I2[54]

  PIN I2[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.144 0.000 64.296 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.144 0.000 64.296 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.144 0.000 64.296 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.144 0.000 64.296 0.152 ;
    END
  END I2[55]

  PIN I2[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.880 0.000 67.032 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.880 0.000 67.032 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.880 0.000 67.032 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.880 0.000 67.032 0.152 ;
    END
  END I2[56]

  PIN I2[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.184 0.000 67.336 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.184 0.000 67.336 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.184 0.000 67.336 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.184 0.000 67.336 0.152 ;
    END
  END I2[57]

  PIN I2[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.488 0.000 67.640 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.488 0.000 67.640 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.488 0.000 67.640 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.488 0.000 67.640 0.152 ;
    END
  END I2[58]

  PIN I2[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.792 0.000 67.944 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.792 0.000 67.944 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.792 0.000 67.944 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.792 0.000 67.944 0.152 ;
    END
  END I2[59]

  PIN I2[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.528 0.000 70.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.528 0.000 70.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.528 0.000 70.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.528 0.000 70.680 0.152 ;
    END
  END I2[60]

  PIN I2[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.832 0.000 70.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.832 0.000 70.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.832 0.000 70.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.832 0.000 70.984 0.152 ;
    END
  END I2[61]

  PIN I2[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.136 0.000 71.288 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.136 0.000 71.288 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.136 0.000 71.288 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.136 0.000 71.288 0.152 ;
    END
  END I2[62]

  PIN I2[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.440 0.000 71.592 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.440 0.000 71.592 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.440 0.000 71.592 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.440 0.000 71.592 0.152 ;
    END
  END I2[63]

  PIN I2[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.176 0.000 74.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.176 0.000 74.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.176 0.000 74.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.176 0.000 74.328 0.152 ;
    END
  END I2[64]

  PIN I2[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.480 0.000 74.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.480 0.000 74.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.480 0.000 74.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.480 0.000 74.632 0.152 ;
    END
  END I2[65]

  PIN I2[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.784 0.000 74.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.784 0.000 74.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.784 0.000 74.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.784 0.000 74.936 0.152 ;
    END
  END I2[66]

  PIN I2[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.088 0.000 75.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 75.088 0.000 75.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 75.088 0.000 75.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 75.088 0.000 75.240 0.152 ;
    END
  END I2[67]

  PIN I2[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.824 0.000 77.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.824 0.000 77.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.824 0.000 77.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.824 0.000 77.976 0.152 ;
    END
  END I2[68]

  PIN I2[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.128 0.000 78.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.128 0.000 78.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.128 0.000 78.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.128 0.000 78.280 0.152 ;
    END
  END I2[69]

  PIN I2[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.432 0.000 78.584 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.432 0.000 78.584 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.432 0.000 78.584 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.432 0.000 78.584 0.152 ;
    END
  END I2[70]

  PIN I2[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.736 0.000 78.888 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.736 0.000 78.888 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.736 0.000 78.888 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.736 0.000 78.888 0.152 ;
    END
  END I2[71]

  PIN I2[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.472 0.000 81.624 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.472 0.000 81.624 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.472 0.000 81.624 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.472 0.000 81.624 0.152 ;
    END
  END I2[72]

  PIN I2[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.776 0.000 81.928 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.776 0.000 81.928 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.776 0.000 81.928 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.776 0.000 81.928 0.152 ;
    END
  END I2[73]

  PIN I2[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.080 0.000 82.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.080 0.000 82.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.080 0.000 82.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.080 0.000 82.232 0.152 ;
    END
  END I2[74]

  PIN I2[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
  END I2[75]

  PIN I2[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.120 0.000 85.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.120 0.000 85.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.120 0.000 85.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.120 0.000 85.272 0.152 ;
    END
  END I2[76]

  PIN I2[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.424 0.000 85.576 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.424 0.000 85.576 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.424 0.000 85.576 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.424 0.000 85.576 0.152 ;
    END
  END I2[77]

  PIN I2[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.728 0.000 85.880 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.728 0.000 85.880 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.728 0.000 85.880 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.728 0.000 85.880 0.152 ;
    END
  END I2[78]

  PIN I2[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.032 0.000 86.184 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.032 0.000 86.184 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.032 0.000 86.184 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.032 0.000 86.184 0.152 ;
    END
  END I2[79]

  PIN I2[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
  END I2[80]

  PIN I2[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.072 0.000 89.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.072 0.000 89.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.072 0.000 89.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.072 0.000 89.224 0.152 ;
    END
  END I2[81]

  PIN I2[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.376 0.000 89.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.376 0.000 89.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.376 0.000 89.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.376 0.000 89.528 0.152 ;
    END
  END I2[82]

  PIN I2[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.680 0.000 89.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.680 0.000 89.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.680 0.000 89.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.680 0.000 89.832 0.152 ;
    END
  END I2[83]

  PIN I2[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.416 0.000 92.568 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.416 0.000 92.568 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.416 0.000 92.568 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.416 0.000 92.568 0.152 ;
    END
  END I2[84]

  PIN I2[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 92.720 0.000 92.872 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 92.720 0.000 92.872 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 92.720 0.000 92.872 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 92.720 0.000 92.872 0.152 ;
    END
  END I2[85]

  PIN I2[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
  END I2[86]

  PIN I2[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.328 0.000 93.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.328 0.000 93.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.328 0.000 93.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.328 0.000 93.480 0.152 ;
    END
  END I2[87]

  PIN I2[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.064 0.000 96.216 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.064 0.000 96.216 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.064 0.000 96.216 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.064 0.000 96.216 0.152 ;
    END
  END I2[88]

  PIN I2[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.368 0.000 96.520 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.368 0.000 96.520 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.368 0.000 96.520 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.368 0.000 96.520 0.152 ;
    END
  END I2[89]

  PIN I2[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.672 0.000 96.824 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.672 0.000 96.824 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.672 0.000 96.824 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.672 0.000 96.824 0.152 ;
    END
  END I2[90]

  PIN I2[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.976 0.000 97.128 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.976 0.000 97.128 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.976 0.000 97.128 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.976 0.000 97.128 0.152 ;
    END
  END I2[91]

  PIN I2[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.712 0.000 99.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.712 0.000 99.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.712 0.000 99.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.712 0.000 99.864 0.152 ;
    END
  END I2[92]

  PIN I2[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.016 0.000 100.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.016 0.000 100.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.016 0.000 100.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.016 0.000 100.168 0.152 ;
    END
  END I2[93]

  PIN I2[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.320 0.000 100.472 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.320 0.000 100.472 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.320 0.000 100.472 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.320 0.000 100.472 0.152 ;
    END
  END I2[94]

  PIN I2[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.624 0.000 100.776 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.624 0.000 100.776 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.624 0.000 100.776 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.624 0.000 100.776 0.152 ;
    END
  END I2[95]

  PIN I2[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.360 0.000 103.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.360 0.000 103.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.360 0.000 103.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.360 0.000 103.512 0.152 ;
    END
  END I2[96]

  PIN I2[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.664 0.000 103.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.664 0.000 103.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.664 0.000 103.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.664 0.000 103.816 0.152 ;
    END
  END I2[97]

  PIN I2[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.968 0.000 104.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.968 0.000 104.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.968 0.000 104.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.968 0.000 104.120 0.152 ;
    END
  END I2[98]

  PIN I2[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.272 0.000 104.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.272 0.000 104.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.272 0.000 104.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.272 0.000 104.424 0.152 ;
    END
  END I2[99]

  PIN I2[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.008 0.000 107.160 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.008 0.000 107.160 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.008 0.000 107.160 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.008 0.000 107.160 0.152 ;
    END
  END I2[100]

  PIN I2[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.312 0.000 107.464 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.312 0.000 107.464 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.312 0.000 107.464 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.312 0.000 107.464 0.152 ;
    END
  END I2[101]

  PIN I2[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.616 0.000 107.768 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.616 0.000 107.768 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.616 0.000 107.768 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.616 0.000 107.768 0.152 ;
    END
  END I2[102]

  PIN I2[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.920 0.000 108.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.920 0.000 108.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.920 0.000 108.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.920 0.000 108.072 0.152 ;
    END
  END I2[103]

  PIN I2[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.656 0.000 110.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.656 0.000 110.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.656 0.000 110.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.656 0.000 110.808 0.152 ;
    END
  END I2[104]

  PIN I2[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.960 0.000 111.112 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.960 0.000 111.112 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.960 0.000 111.112 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.960 0.000 111.112 0.152 ;
    END
  END I2[105]

  PIN I2[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.264 0.000 111.416 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 111.264 0.000 111.416 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 111.264 0.000 111.416 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.264 0.000 111.416 0.152 ;
    END
  END I2[106]

  PIN I2[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.568 0.000 111.720 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 111.568 0.000 111.720 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 111.568 0.000 111.720 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.568 0.000 111.720 0.152 ;
    END
  END I2[107]

  PIN I2[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.304 0.000 114.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 114.304 0.000 114.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 114.304 0.000 114.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.304 0.000 114.456 0.152 ;
    END
  END I2[108]

  PIN I2[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.608 0.000 114.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 114.608 0.000 114.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 114.608 0.000 114.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.608 0.000 114.760 0.152 ;
    END
  END I2[109]

  PIN I2[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.912 0.000 115.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 114.912 0.000 115.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 114.912 0.000 115.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.912 0.000 115.064 0.152 ;
    END
  END I2[110]

  PIN I2[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.216 0.000 115.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 115.216 0.000 115.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 115.216 0.000 115.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.216 0.000 115.368 0.152 ;
    END
  END I2[111]

  PIN I2[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.952 0.000 118.104 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 117.952 0.000 118.104 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 117.952 0.000 118.104 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.952 0.000 118.104 0.152 ;
    END
  END I2[112]

  PIN I2[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.256 0.000 118.408 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 118.256 0.000 118.408 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 118.256 0.000 118.408 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.256 0.000 118.408 0.152 ;
    END
  END I2[113]

  PIN I2[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.560 0.000 118.712 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 118.560 0.000 118.712 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 118.560 0.000 118.712 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.560 0.000 118.712 0.152 ;
    END
  END I2[114]

  PIN I2[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.864 0.000 119.016 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 118.864 0.000 119.016 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 118.864 0.000 119.016 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.864 0.000 119.016 0.152 ;
    END
  END I2[115]

  PIN I2[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.600 0.000 121.752 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 121.600 0.000 121.752 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 121.600 0.000 121.752 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.600 0.000 121.752 0.152 ;
    END
  END I2[116]

  PIN I2[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.904 0.000 122.056 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 121.904 0.000 122.056 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 121.904 0.000 122.056 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.904 0.000 122.056 0.152 ;
    END
  END I2[117]

  PIN I2[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.208 0.000 122.360 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 122.208 0.000 122.360 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 122.208 0.000 122.360 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.208 0.000 122.360 0.152 ;
    END
  END I2[118]

  PIN I2[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.512 0.000 122.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 122.512 0.000 122.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 122.512 0.000 122.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.512 0.000 122.664 0.152 ;
    END
  END I2[119]

  PIN I2[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.248 0.000 125.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 125.248 0.000 125.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 125.248 0.000 125.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.248 0.000 125.400 0.152 ;
    END
  END I2[120]

  PIN I2[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.552 0.000 125.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 125.552 0.000 125.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 125.552 0.000 125.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.552 0.000 125.704 0.152 ;
    END
  END I2[121]

  PIN I2[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.856 0.000 126.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 125.856 0.000 126.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 125.856 0.000 126.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.856 0.000 126.008 0.152 ;
    END
  END I2[122]

  PIN I2[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.160 0.000 126.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 126.160 0.000 126.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 126.160 0.000 126.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.160 0.000 126.312 0.152 ;
    END
  END I2[123]

  PIN I2[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.896 0.000 129.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 128.896 0.000 129.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 128.896 0.000 129.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 128.896 0.000 129.048 0.152 ;
    END
  END I2[124]

  PIN I2[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.200 0.000 129.352 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 129.200 0.000 129.352 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 129.200 0.000 129.352 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.200 0.000 129.352 0.152 ;
    END
  END I2[125]

  PIN I2[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.504 0.000 129.656 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 129.504 0.000 129.656 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 129.504 0.000 129.656 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.504 0.000 129.656 0.152 ;
    END
  END I2[126]

  PIN I2[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.808 0.000 129.960 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 129.808 0.000 129.960 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 129.808 0.000 129.960 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.808 0.000 129.960 0.152 ;
    END
  END I2[127]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 119.168 0.152 119.320 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 119.168 0.152 119.320 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 119.168 0.152 119.320 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 119.168 0.152 119.320 ;
    END
  END A2[0]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 115.520 0.152 115.672 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 115.520 0.152 115.672 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 115.520 0.152 115.672 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 115.520 0.152 115.672 ;
    END
  END A2[1]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 111.872 0.152 112.024 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 111.872 0.152 112.024 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 111.872 0.152 112.024 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 111.872 0.152 112.024 ;
    END
  END A2[2]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 108.224 0.152 108.376 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 108.224 0.152 108.376 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 108.224 0.152 108.376 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 108.224 0.152 108.376 ;
    END
  END A2[3]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 104.576 0.152 104.728 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 104.576 0.152 104.728 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 104.576 0.152 104.728 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 104.576 0.152 104.728 ;
    END
  END A2[4]

  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 100.928 0.152 101.080 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 100.928 0.152 101.080 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 100.928 0.152 101.080 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 100.928 0.152 101.080 ;
    END
  END A2[5]

  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 97.280 0.152 97.432 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 97.280 0.152 97.432 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 97.280 0.152 97.432 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 97.280 0.152 97.432 ;
    END
  END A2[6]

  PIN A2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 93.632 0.152 93.784 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 93.632 0.152 93.784 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 93.632 0.152 93.784 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 93.632 0.152 93.784 ;
    END
  END A2[7]

  PIN A2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 89.984 0.152 90.136 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 89.984 0.152 90.136 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 89.984 0.152 90.136 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 89.984 0.152 90.136 ;
    END
  END A2[8]

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 34.048 0.152 34.200 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 34.048 0.152 34.200 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 34.048 0.152 34.200 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 34.048 0.152 34.200 ;
    END
  END WEB2

  PIN WBM2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 32.832 0.152 32.984 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 32.832 0.152 32.984 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 32.832 0.152 32.984 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 32.832 0.152 32.984 ;
    END
  END WBM2[0]

  PIN WBM2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 31.616 0.152 31.768 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 31.616 0.152 31.768 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 31.616 0.152 31.768 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 31.616 0.152 31.768 ;
    END
  END WBM2[1]

  PIN WBM2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 30.400 0.152 30.552 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 30.400 0.152 30.552 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 30.400 0.152 30.552 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 30.400 0.152 30.552 ;
    END
  END WBM2[2]

  PIN WBM2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 29.184 0.152 29.336 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 29.184 0.152 29.336 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 29.184 0.152 29.336 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 29.184 0.152 29.336 ;
    END
  END WBM2[3]

  PIN WBM2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 27.968 0.152 28.120 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 27.968 0.152 28.120 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 27.968 0.152 28.120 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 27.968 0.152 28.120 ;
    END
  END WBM2[4]

  PIN WBM2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 26.752 0.152 26.904 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 26.752 0.152 26.904 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 26.752 0.152 26.904 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 26.752 0.152 26.904 ;
    END
  END WBM2[5]

  PIN WBM2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 25.536 0.152 25.688 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 25.536 0.152 25.688 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 25.536 0.152 25.688 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 25.536 0.152 25.688 ;
    END
  END WBM2[6]

  PIN WBM2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 24.320 0.152 24.472 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 24.320 0.152 24.472 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 24.320 0.152 24.472 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 24.320 0.152 24.472 ;
    END
  END WBM2[7]

  PIN WBM2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 23.104 0.152 23.256 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 23.104 0.152 23.256 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 23.104 0.152 23.256 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 23.104 0.152 23.256 ;
    END
  END WBM2[8]

  PIN WBM2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 21.888 0.152 22.040 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 21.888 0.152 22.040 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 21.888 0.152 22.040 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 21.888 0.152 22.040 ;
    END
  END WBM2[9]

  PIN WBM2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 20.672 0.152 20.824 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 20.672 0.152 20.824 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 20.672 0.152 20.824 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 20.672 0.152 20.824 ;
    END
  END WBM2[10]

  PIN WBM2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 19.456 0.152 19.608 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 19.456 0.152 19.608 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 19.456 0.152 19.608 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 19.456 0.152 19.608 ;
    END
  END WBM2[11]

  PIN WBM2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 18.240 0.152 18.392 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 18.240 0.152 18.392 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 18.240 0.152 18.392 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 18.240 0.152 18.392 ;
    END
  END WBM2[12]

  PIN WBM2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 17.024 0.152 17.176 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 17.024 0.152 17.176 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 17.024 0.152 17.176 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 17.024 0.152 17.176 ;
    END
  END WBM2[13]

  PIN WBM2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 15.808 0.152 15.960 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 15.808 0.152 15.960 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 15.808 0.152 15.960 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 15.808 0.152 15.960 ;
    END
  END WBM2[14]

  PIN WBM2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 14.592 0.152 14.744 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 14.592 0.152 14.744 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 14.592 0.152 14.744 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 14.592 0.152 14.744 ;
    END
  END WBM2[15]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 5.195 134.192 7.195 136.192 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.195 134.192 7.195 136.192 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.195 134.192 7.195 136.192 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M2 ;
        RECT 7.915 134.192 9.915 136.192 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.915 134.192 9.915 136.192 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.915 134.192 9.915 136.192 ;
    END
  END VSS

  OBS
    LAYER M2 ;
      RECT 268.432 0.000 278.464 0.304 ;
      RECT 265.696 0.000 267.976 0.304 ;
      RECT 262.960 0.000 265.240 0.304 ;
      RECT 260.224 0.000 262.504 0.304 ;
      RECT 256.576 0.000 258.856 0.304 ;
      RECT 252.928 0.000 255.208 0.304 ;
      RECT 249.280 0.000 251.560 0.304 ;
      RECT 245.632 0.000 247.912 0.304 ;
      RECT 241.984 0.000 244.264 0.304 ;
      RECT 238.336 0.000 240.616 0.304 ;
      RECT 234.688 0.000 236.968 0.304 ;
      RECT 231.040 0.000 233.320 0.304 ;
      RECT 227.392 0.000 229.672 0.304 ;
      RECT 223.744 0.000 226.024 0.304 ;
      RECT 220.096 0.000 222.376 0.304 ;
      RECT 216.448 0.000 218.728 0.304 ;
      RECT 212.800 0.000 215.080 0.304 ;
      RECT 209.152 0.000 211.432 0.304 ;
      RECT 205.504 0.000 207.784 0.304 ;
      RECT 201.856 0.000 204.136 0.304 ;
      RECT 198.208 0.000 200.488 0.304 ;
      RECT 194.560 0.000 196.840 0.304 ;
      RECT 190.912 0.000 193.192 0.304 ;
      RECT 187.264 0.000 189.544 0.304 ;
      RECT 183.616 0.000 185.896 0.304 ;
      RECT 179.968 0.000 182.248 0.304 ;
      RECT 176.320 0.000 178.600 0.304 ;
      RECT 172.672 0.000 174.952 0.304 ;
      RECT 169.024 0.000 171.304 0.304 ;
      RECT 165.376 0.000 167.656 0.304 ;
      RECT 161.728 0.000 164.008 0.304 ;
      RECT 158.080 0.000 160.360 0.304 ;
      RECT 154.432 0.000 156.712 0.304 ;
      RECT 150.784 0.000 153.064 0.304 ;
      RECT 147.136 0.000 149.416 0.304 ;
      RECT 278.160 119.472 278.464 134.040 ;
      RECT 278.160 115.824 278.464 119.016 ;
      RECT 278.160 112.176 278.464 115.368 ;
      RECT 278.160 108.528 278.464 111.720 ;
      RECT 278.160 104.880 278.464 108.072 ;
      RECT 278.160 101.232 278.464 104.424 ;
      RECT 278.160 97.584 278.464 100.776 ;
      RECT 278.160 93.936 278.464 97.128 ;
      RECT 278.160 90.288 278.464 93.480 ;
      RECT 278.160 34.352 278.464 89.832 ;
      RECT 278.160 33.136 278.464 33.896 ;
      RECT 278.160 31.920 278.464 32.680 ;
      RECT 278.160 30.704 278.464 31.464 ;
      RECT 278.160 29.488 278.464 30.248 ;
      RECT 278.160 28.272 278.464 29.032 ;
      RECT 278.160 27.056 278.464 27.816 ;
      RECT 278.160 25.840 278.464 26.600 ;
      RECT 278.160 24.624 278.464 25.384 ;
      RECT 278.160 23.408 278.464 24.168 ;
      RECT 278.160 22.192 278.464 22.952 ;
      RECT 278.160 20.976 278.464 21.736 ;
      RECT 278.160 19.760 278.464 20.520 ;
      RECT 278.160 18.544 278.464 19.304 ;
      RECT 278.160 17.328 278.464 18.088 ;
      RECT 278.160 16.112 278.464 16.872 ;
      RECT 278.160 14.896 278.464 15.656 ;
      RECT 278.160 0.304 278.464 14.440 ;
      RECT 0.000 0.000 10.184 0.304 ;
      RECT 10.640 0.000 12.920 0.304 ;
      RECT 13.376 0.000 15.656 0.304 ;
      RECT 17.024 0.000 19.304 0.304 ;
      RECT 20.672 0.000 22.952 0.304 ;
      RECT 24.320 0.000 26.600 0.304 ;
      RECT 27.968 0.000 30.248 0.304 ;
      RECT 31.616 0.000 33.896 0.304 ;
      RECT 35.264 0.000 37.544 0.304 ;
      RECT 38.912 0.000 41.192 0.304 ;
      RECT 42.560 0.000 44.840 0.304 ;
      RECT 46.208 0.000 48.488 0.304 ;
      RECT 49.856 0.000 52.136 0.304 ;
      RECT 53.504 0.000 55.784 0.304 ;
      RECT 57.152 0.000 59.432 0.304 ;
      RECT 60.800 0.000 63.080 0.304 ;
      RECT 64.448 0.000 66.728 0.304 ;
      RECT 68.096 0.000 70.376 0.304 ;
      RECT 71.744 0.000 74.024 0.304 ;
      RECT 75.392 0.000 77.672 0.304 ;
      RECT 79.040 0.000 81.320 0.304 ;
      RECT 82.688 0.000 84.968 0.304 ;
      RECT 86.336 0.000 88.616 0.304 ;
      RECT 89.984 0.000 92.264 0.304 ;
      RECT 93.632 0.000 95.912 0.304 ;
      RECT 97.280 0.000 99.560 0.304 ;
      RECT 100.928 0.000 103.208 0.304 ;
      RECT 104.576 0.000 106.856 0.304 ;
      RECT 108.224 0.000 110.504 0.304 ;
      RECT 111.872 0.000 114.152 0.304 ;
      RECT 115.520 0.000 117.800 0.304 ;
      RECT 119.168 0.000 121.448 0.304 ;
      RECT 122.816 0.000 125.096 0.304 ;
      RECT 126.464 0.000 128.744 0.304 ;
      RECT 130.112 0.000 145.768 0.304 ;
      RECT 0.000 119.472 0.304 134.040 ;
      RECT 0.000 115.824 0.304 119.016 ;
      RECT 0.000 112.176 0.304 115.368 ;
      RECT 0.000 108.528 0.304 111.720 ;
      RECT 0.000 104.880 0.304 108.072 ;
      RECT 0.000 101.232 0.304 104.424 ;
      RECT 0.000 97.584 0.304 100.776 ;
      RECT 0.000 93.936 0.304 97.128 ;
      RECT 0.000 90.288 0.304 93.480 ;
      RECT 0.000 34.352 0.304 89.832 ;
      RECT 0.000 33.136 0.304 33.896 ;
      RECT 0.000 31.920 0.304 32.680 ;
      RECT 0.000 30.704 0.304 31.464 ;
      RECT 0.000 29.488 0.304 30.248 ;
      RECT 0.000 28.272 0.304 29.032 ;
      RECT 0.000 27.056 0.304 27.816 ;
      RECT 0.000 25.840 0.304 26.600 ;
      RECT 0.000 24.624 0.304 25.384 ;
      RECT 0.000 23.408 0.304 24.168 ;
      RECT 0.000 22.192 0.304 22.952 ;
      RECT 0.000 20.976 0.304 21.736 ;
      RECT 0.000 19.760 0.304 20.520 ;
      RECT 0.000 18.544 0.304 19.304 ;
      RECT 0.000 17.328 0.304 18.088 ;
      RECT 0.000 16.112 0.304 16.872 ;
      RECT 0.000 14.896 0.304 15.656 ;
      RECT 0.000 0.304 0.304 14.440 ;
      RECT 0.000 134.040 5.043 136.192 ;
      RECT 7.355 134.040 7.763 136.192 ;
      RECT 10.067 134.040 278.464 136.192 ;
      RECT 0.304 0.304 278.160 134.040 ;
    LAYER M3 ;
      RECT 268.432 0.000 278.464 0.304 ;
      RECT 265.696 0.000 267.976 0.304 ;
      RECT 262.960 0.000 265.240 0.304 ;
      RECT 260.224 0.000 262.504 0.304 ;
      RECT 256.576 0.000 258.856 0.304 ;
      RECT 252.928 0.000 255.208 0.304 ;
      RECT 249.280 0.000 251.560 0.304 ;
      RECT 245.632 0.000 247.912 0.304 ;
      RECT 241.984 0.000 244.264 0.304 ;
      RECT 238.336 0.000 240.616 0.304 ;
      RECT 234.688 0.000 236.968 0.304 ;
      RECT 231.040 0.000 233.320 0.304 ;
      RECT 227.392 0.000 229.672 0.304 ;
      RECT 223.744 0.000 226.024 0.304 ;
      RECT 220.096 0.000 222.376 0.304 ;
      RECT 216.448 0.000 218.728 0.304 ;
      RECT 212.800 0.000 215.080 0.304 ;
      RECT 209.152 0.000 211.432 0.304 ;
      RECT 205.504 0.000 207.784 0.304 ;
      RECT 201.856 0.000 204.136 0.304 ;
      RECT 198.208 0.000 200.488 0.304 ;
      RECT 194.560 0.000 196.840 0.304 ;
      RECT 190.912 0.000 193.192 0.304 ;
      RECT 187.264 0.000 189.544 0.304 ;
      RECT 183.616 0.000 185.896 0.304 ;
      RECT 179.968 0.000 182.248 0.304 ;
      RECT 176.320 0.000 178.600 0.304 ;
      RECT 172.672 0.000 174.952 0.304 ;
      RECT 169.024 0.000 171.304 0.304 ;
      RECT 165.376 0.000 167.656 0.304 ;
      RECT 161.728 0.000 164.008 0.304 ;
      RECT 158.080 0.000 160.360 0.304 ;
      RECT 154.432 0.000 156.712 0.304 ;
      RECT 150.784 0.000 153.064 0.304 ;
      RECT 147.136 0.000 149.416 0.304 ;
      RECT 278.160 119.472 278.464 134.040 ;
      RECT 278.160 115.824 278.464 119.016 ;
      RECT 278.160 112.176 278.464 115.368 ;
      RECT 278.160 108.528 278.464 111.720 ;
      RECT 278.160 104.880 278.464 108.072 ;
      RECT 278.160 101.232 278.464 104.424 ;
      RECT 278.160 97.584 278.464 100.776 ;
      RECT 278.160 93.936 278.464 97.128 ;
      RECT 278.160 90.288 278.464 93.480 ;
      RECT 278.160 34.352 278.464 89.832 ;
      RECT 278.160 33.136 278.464 33.896 ;
      RECT 278.160 31.920 278.464 32.680 ;
      RECT 278.160 30.704 278.464 31.464 ;
      RECT 278.160 29.488 278.464 30.248 ;
      RECT 278.160 28.272 278.464 29.032 ;
      RECT 278.160 27.056 278.464 27.816 ;
      RECT 278.160 25.840 278.464 26.600 ;
      RECT 278.160 24.624 278.464 25.384 ;
      RECT 278.160 23.408 278.464 24.168 ;
      RECT 278.160 22.192 278.464 22.952 ;
      RECT 278.160 20.976 278.464 21.736 ;
      RECT 278.160 19.760 278.464 20.520 ;
      RECT 278.160 18.544 278.464 19.304 ;
      RECT 278.160 17.328 278.464 18.088 ;
      RECT 278.160 16.112 278.464 16.872 ;
      RECT 278.160 14.896 278.464 15.656 ;
      RECT 278.160 0.304 278.464 14.440 ;
      RECT 0.000 0.000 10.184 0.304 ;
      RECT 10.640 0.000 12.920 0.304 ;
      RECT 13.376 0.000 15.656 0.304 ;
      RECT 17.024 0.000 19.304 0.304 ;
      RECT 20.672 0.000 22.952 0.304 ;
      RECT 24.320 0.000 26.600 0.304 ;
      RECT 27.968 0.000 30.248 0.304 ;
      RECT 31.616 0.000 33.896 0.304 ;
      RECT 35.264 0.000 37.544 0.304 ;
      RECT 38.912 0.000 41.192 0.304 ;
      RECT 42.560 0.000 44.840 0.304 ;
      RECT 46.208 0.000 48.488 0.304 ;
      RECT 49.856 0.000 52.136 0.304 ;
      RECT 53.504 0.000 55.784 0.304 ;
      RECT 57.152 0.000 59.432 0.304 ;
      RECT 60.800 0.000 63.080 0.304 ;
      RECT 64.448 0.000 66.728 0.304 ;
      RECT 68.096 0.000 70.376 0.304 ;
      RECT 71.744 0.000 74.024 0.304 ;
      RECT 75.392 0.000 77.672 0.304 ;
      RECT 79.040 0.000 81.320 0.304 ;
      RECT 82.688 0.000 84.968 0.304 ;
      RECT 86.336 0.000 88.616 0.304 ;
      RECT 89.984 0.000 92.264 0.304 ;
      RECT 93.632 0.000 95.912 0.304 ;
      RECT 97.280 0.000 99.560 0.304 ;
      RECT 100.928 0.000 103.208 0.304 ;
      RECT 104.576 0.000 106.856 0.304 ;
      RECT 108.224 0.000 110.504 0.304 ;
      RECT 111.872 0.000 114.152 0.304 ;
      RECT 115.520 0.000 117.800 0.304 ;
      RECT 119.168 0.000 121.448 0.304 ;
      RECT 122.816 0.000 125.096 0.304 ;
      RECT 126.464 0.000 128.744 0.304 ;
      RECT 130.112 0.000 145.768 0.304 ;
      RECT 0.000 119.472 0.304 134.040 ;
      RECT 0.000 115.824 0.304 119.016 ;
      RECT 0.000 112.176 0.304 115.368 ;
      RECT 0.000 108.528 0.304 111.720 ;
      RECT 0.000 104.880 0.304 108.072 ;
      RECT 0.000 101.232 0.304 104.424 ;
      RECT 0.000 97.584 0.304 100.776 ;
      RECT 0.000 93.936 0.304 97.128 ;
      RECT 0.000 90.288 0.304 93.480 ;
      RECT 0.000 34.352 0.304 89.832 ;
      RECT 0.000 33.136 0.304 33.896 ;
      RECT 0.000 31.920 0.304 32.680 ;
      RECT 0.000 30.704 0.304 31.464 ;
      RECT 0.000 29.488 0.304 30.248 ;
      RECT 0.000 28.272 0.304 29.032 ;
      RECT 0.000 27.056 0.304 27.816 ;
      RECT 0.000 25.840 0.304 26.600 ;
      RECT 0.000 24.624 0.304 25.384 ;
      RECT 0.000 23.408 0.304 24.168 ;
      RECT 0.000 22.192 0.304 22.952 ;
      RECT 0.000 20.976 0.304 21.736 ;
      RECT 0.000 19.760 0.304 20.520 ;
      RECT 0.000 18.544 0.304 19.304 ;
      RECT 0.000 17.328 0.304 18.088 ;
      RECT 0.000 16.112 0.304 16.872 ;
      RECT 0.000 14.896 0.304 15.656 ;
      RECT 0.000 0.304 0.304 14.440 ;
      RECT 0.000 134.040 5.043 136.192 ;
      RECT 7.355 134.040 7.763 136.192 ;
      RECT 10.067 134.040 278.464 136.192 ;
      RECT 0.304 0.304 278.160 134.040 ;
    LAYER M4 ;
      RECT 268.432 0.000 278.464 0.304 ;
      RECT 265.696 0.000 267.976 0.304 ;
      RECT 262.960 0.000 265.240 0.304 ;
      RECT 260.224 0.000 262.504 0.304 ;
      RECT 256.576 0.000 258.856 0.304 ;
      RECT 252.928 0.000 255.208 0.304 ;
      RECT 249.280 0.000 251.560 0.304 ;
      RECT 245.632 0.000 247.912 0.304 ;
      RECT 241.984 0.000 244.264 0.304 ;
      RECT 238.336 0.000 240.616 0.304 ;
      RECT 234.688 0.000 236.968 0.304 ;
      RECT 231.040 0.000 233.320 0.304 ;
      RECT 227.392 0.000 229.672 0.304 ;
      RECT 223.744 0.000 226.024 0.304 ;
      RECT 220.096 0.000 222.376 0.304 ;
      RECT 216.448 0.000 218.728 0.304 ;
      RECT 212.800 0.000 215.080 0.304 ;
      RECT 209.152 0.000 211.432 0.304 ;
      RECT 205.504 0.000 207.784 0.304 ;
      RECT 201.856 0.000 204.136 0.304 ;
      RECT 198.208 0.000 200.488 0.304 ;
      RECT 194.560 0.000 196.840 0.304 ;
      RECT 190.912 0.000 193.192 0.304 ;
      RECT 187.264 0.000 189.544 0.304 ;
      RECT 183.616 0.000 185.896 0.304 ;
      RECT 179.968 0.000 182.248 0.304 ;
      RECT 176.320 0.000 178.600 0.304 ;
      RECT 172.672 0.000 174.952 0.304 ;
      RECT 169.024 0.000 171.304 0.304 ;
      RECT 165.376 0.000 167.656 0.304 ;
      RECT 161.728 0.000 164.008 0.304 ;
      RECT 158.080 0.000 160.360 0.304 ;
      RECT 154.432 0.000 156.712 0.304 ;
      RECT 150.784 0.000 153.064 0.304 ;
      RECT 147.136 0.000 149.416 0.304 ;
      RECT 278.160 119.472 278.464 134.040 ;
      RECT 278.160 115.824 278.464 119.016 ;
      RECT 278.160 112.176 278.464 115.368 ;
      RECT 278.160 108.528 278.464 111.720 ;
      RECT 278.160 104.880 278.464 108.072 ;
      RECT 278.160 101.232 278.464 104.424 ;
      RECT 278.160 97.584 278.464 100.776 ;
      RECT 278.160 93.936 278.464 97.128 ;
      RECT 278.160 90.288 278.464 93.480 ;
      RECT 278.160 34.352 278.464 89.832 ;
      RECT 278.160 33.136 278.464 33.896 ;
      RECT 278.160 31.920 278.464 32.680 ;
      RECT 278.160 30.704 278.464 31.464 ;
      RECT 278.160 29.488 278.464 30.248 ;
      RECT 278.160 28.272 278.464 29.032 ;
      RECT 278.160 27.056 278.464 27.816 ;
      RECT 278.160 25.840 278.464 26.600 ;
      RECT 278.160 24.624 278.464 25.384 ;
      RECT 278.160 23.408 278.464 24.168 ;
      RECT 278.160 22.192 278.464 22.952 ;
      RECT 278.160 20.976 278.464 21.736 ;
      RECT 278.160 19.760 278.464 20.520 ;
      RECT 278.160 18.544 278.464 19.304 ;
      RECT 278.160 17.328 278.464 18.088 ;
      RECT 278.160 16.112 278.464 16.872 ;
      RECT 278.160 14.896 278.464 15.656 ;
      RECT 278.160 0.304 278.464 14.440 ;
      RECT 0.000 0.000 10.184 0.304 ;
      RECT 10.640 0.000 12.920 0.304 ;
      RECT 13.376 0.000 15.656 0.304 ;
      RECT 17.024 0.000 19.304 0.304 ;
      RECT 20.672 0.000 22.952 0.304 ;
      RECT 24.320 0.000 26.600 0.304 ;
      RECT 27.968 0.000 30.248 0.304 ;
      RECT 31.616 0.000 33.896 0.304 ;
      RECT 35.264 0.000 37.544 0.304 ;
      RECT 38.912 0.000 41.192 0.304 ;
      RECT 42.560 0.000 44.840 0.304 ;
      RECT 46.208 0.000 48.488 0.304 ;
      RECT 49.856 0.000 52.136 0.304 ;
      RECT 53.504 0.000 55.784 0.304 ;
      RECT 57.152 0.000 59.432 0.304 ;
      RECT 60.800 0.000 63.080 0.304 ;
      RECT 64.448 0.000 66.728 0.304 ;
      RECT 68.096 0.000 70.376 0.304 ;
      RECT 71.744 0.000 74.024 0.304 ;
      RECT 75.392 0.000 77.672 0.304 ;
      RECT 79.040 0.000 81.320 0.304 ;
      RECT 82.688 0.000 84.968 0.304 ;
      RECT 86.336 0.000 88.616 0.304 ;
      RECT 89.984 0.000 92.264 0.304 ;
      RECT 93.632 0.000 95.912 0.304 ;
      RECT 97.280 0.000 99.560 0.304 ;
      RECT 100.928 0.000 103.208 0.304 ;
      RECT 104.576 0.000 106.856 0.304 ;
      RECT 108.224 0.000 110.504 0.304 ;
      RECT 111.872 0.000 114.152 0.304 ;
      RECT 115.520 0.000 117.800 0.304 ;
      RECT 119.168 0.000 121.448 0.304 ;
      RECT 122.816 0.000 125.096 0.304 ;
      RECT 126.464 0.000 128.744 0.304 ;
      RECT 130.112 0.000 145.768 0.304 ;
      RECT 0.000 119.472 0.304 134.040 ;
      RECT 0.000 115.824 0.304 119.016 ;
      RECT 0.000 112.176 0.304 115.368 ;
      RECT 0.000 108.528 0.304 111.720 ;
      RECT 0.000 104.880 0.304 108.072 ;
      RECT 0.000 101.232 0.304 104.424 ;
      RECT 0.000 97.584 0.304 100.776 ;
      RECT 0.000 93.936 0.304 97.128 ;
      RECT 0.000 90.288 0.304 93.480 ;
      RECT 0.000 34.352 0.304 89.832 ;
      RECT 0.000 33.136 0.304 33.896 ;
      RECT 0.000 31.920 0.304 32.680 ;
      RECT 0.000 30.704 0.304 31.464 ;
      RECT 0.000 29.488 0.304 30.248 ;
      RECT 0.000 28.272 0.304 29.032 ;
      RECT 0.000 27.056 0.304 27.816 ;
      RECT 0.000 25.840 0.304 26.600 ;
      RECT 0.000 24.624 0.304 25.384 ;
      RECT 0.000 23.408 0.304 24.168 ;
      RECT 0.000 22.192 0.304 22.952 ;
      RECT 0.000 20.976 0.304 21.736 ;
      RECT 0.000 19.760 0.304 20.520 ;
      RECT 0.000 18.544 0.304 19.304 ;
      RECT 0.000 17.328 0.304 18.088 ;
      RECT 0.000 16.112 0.304 16.872 ;
      RECT 0.000 14.896 0.304 15.656 ;
      RECT 0.000 0.304 0.304 14.440 ;
      RECT 0.000 134.040 5.043 136.192 ;
      RECT 7.355 134.040 7.763 136.192 ;
      RECT 10.067 134.040 278.464 136.192 ;
      RECT 0.304 0.304 278.160 134.040 ;
    LAYER M5 ;
      RECT 268.432 0.000 278.464 0.304 ;
      RECT 265.696 0.000 267.976 0.304 ;
      RECT 262.960 0.000 265.240 0.304 ;
      RECT 260.224 0.000 262.504 0.304 ;
      RECT 256.576 0.000 258.856 0.304 ;
      RECT 252.928 0.000 255.208 0.304 ;
      RECT 249.280 0.000 251.560 0.304 ;
      RECT 245.632 0.000 247.912 0.304 ;
      RECT 241.984 0.000 244.264 0.304 ;
      RECT 238.336 0.000 240.616 0.304 ;
      RECT 234.688 0.000 236.968 0.304 ;
      RECT 231.040 0.000 233.320 0.304 ;
      RECT 227.392 0.000 229.672 0.304 ;
      RECT 223.744 0.000 226.024 0.304 ;
      RECT 220.096 0.000 222.376 0.304 ;
      RECT 216.448 0.000 218.728 0.304 ;
      RECT 212.800 0.000 215.080 0.304 ;
      RECT 209.152 0.000 211.432 0.304 ;
      RECT 205.504 0.000 207.784 0.304 ;
      RECT 201.856 0.000 204.136 0.304 ;
      RECT 198.208 0.000 200.488 0.304 ;
      RECT 194.560 0.000 196.840 0.304 ;
      RECT 190.912 0.000 193.192 0.304 ;
      RECT 187.264 0.000 189.544 0.304 ;
      RECT 183.616 0.000 185.896 0.304 ;
      RECT 179.968 0.000 182.248 0.304 ;
      RECT 176.320 0.000 178.600 0.304 ;
      RECT 172.672 0.000 174.952 0.304 ;
      RECT 169.024 0.000 171.304 0.304 ;
      RECT 165.376 0.000 167.656 0.304 ;
      RECT 161.728 0.000 164.008 0.304 ;
      RECT 158.080 0.000 160.360 0.304 ;
      RECT 154.432 0.000 156.712 0.304 ;
      RECT 150.784 0.000 153.064 0.304 ;
      RECT 147.136 0.000 149.416 0.304 ;
      RECT 278.160 119.472 278.464 134.040 ;
      RECT 278.160 115.824 278.464 119.016 ;
      RECT 278.160 112.176 278.464 115.368 ;
      RECT 278.160 108.528 278.464 111.720 ;
      RECT 278.160 104.880 278.464 108.072 ;
      RECT 278.160 101.232 278.464 104.424 ;
      RECT 278.160 97.584 278.464 100.776 ;
      RECT 278.160 93.936 278.464 97.128 ;
      RECT 278.160 90.288 278.464 93.480 ;
      RECT 278.160 34.352 278.464 89.832 ;
      RECT 278.160 33.136 278.464 33.896 ;
      RECT 278.160 31.920 278.464 32.680 ;
      RECT 278.160 30.704 278.464 31.464 ;
      RECT 278.160 29.488 278.464 30.248 ;
      RECT 278.160 28.272 278.464 29.032 ;
      RECT 278.160 27.056 278.464 27.816 ;
      RECT 278.160 25.840 278.464 26.600 ;
      RECT 278.160 24.624 278.464 25.384 ;
      RECT 278.160 23.408 278.464 24.168 ;
      RECT 278.160 22.192 278.464 22.952 ;
      RECT 278.160 20.976 278.464 21.736 ;
      RECT 278.160 19.760 278.464 20.520 ;
      RECT 278.160 18.544 278.464 19.304 ;
      RECT 278.160 17.328 278.464 18.088 ;
      RECT 278.160 16.112 278.464 16.872 ;
      RECT 278.160 14.896 278.464 15.656 ;
      RECT 278.160 0.304 278.464 14.440 ;
      RECT 0.000 0.000 10.184 0.304 ;
      RECT 10.640 0.000 12.920 0.304 ;
      RECT 13.376 0.000 15.656 0.304 ;
      RECT 17.024 0.000 19.304 0.304 ;
      RECT 20.672 0.000 22.952 0.304 ;
      RECT 24.320 0.000 26.600 0.304 ;
      RECT 27.968 0.000 30.248 0.304 ;
      RECT 31.616 0.000 33.896 0.304 ;
      RECT 35.264 0.000 37.544 0.304 ;
      RECT 38.912 0.000 41.192 0.304 ;
      RECT 42.560 0.000 44.840 0.304 ;
      RECT 46.208 0.000 48.488 0.304 ;
      RECT 49.856 0.000 52.136 0.304 ;
      RECT 53.504 0.000 55.784 0.304 ;
      RECT 57.152 0.000 59.432 0.304 ;
      RECT 60.800 0.000 63.080 0.304 ;
      RECT 64.448 0.000 66.728 0.304 ;
      RECT 68.096 0.000 70.376 0.304 ;
      RECT 71.744 0.000 74.024 0.304 ;
      RECT 75.392 0.000 77.672 0.304 ;
      RECT 79.040 0.000 81.320 0.304 ;
      RECT 82.688 0.000 84.968 0.304 ;
      RECT 86.336 0.000 88.616 0.304 ;
      RECT 89.984 0.000 92.264 0.304 ;
      RECT 93.632 0.000 95.912 0.304 ;
      RECT 97.280 0.000 99.560 0.304 ;
      RECT 100.928 0.000 103.208 0.304 ;
      RECT 104.576 0.000 106.856 0.304 ;
      RECT 108.224 0.000 110.504 0.304 ;
      RECT 111.872 0.000 114.152 0.304 ;
      RECT 115.520 0.000 117.800 0.304 ;
      RECT 119.168 0.000 121.448 0.304 ;
      RECT 122.816 0.000 125.096 0.304 ;
      RECT 126.464 0.000 128.744 0.304 ;
      RECT 130.112 0.000 145.768 0.304 ;
      RECT 0.000 119.472 0.304 134.040 ;
      RECT 0.000 115.824 0.304 119.016 ;
      RECT 0.000 112.176 0.304 115.368 ;
      RECT 0.000 108.528 0.304 111.720 ;
      RECT 0.000 104.880 0.304 108.072 ;
      RECT 0.000 101.232 0.304 104.424 ;
      RECT 0.000 97.584 0.304 100.776 ;
      RECT 0.000 93.936 0.304 97.128 ;
      RECT 0.000 90.288 0.304 93.480 ;
      RECT 0.000 34.352 0.304 89.832 ;
      RECT 0.000 33.136 0.304 33.896 ;
      RECT 0.000 31.920 0.304 32.680 ;
      RECT 0.000 30.704 0.304 31.464 ;
      RECT 0.000 29.488 0.304 30.248 ;
      RECT 0.000 28.272 0.304 29.032 ;
      RECT 0.000 27.056 0.304 27.816 ;
      RECT 0.000 25.840 0.304 26.600 ;
      RECT 0.000 24.624 0.304 25.384 ;
      RECT 0.000 23.408 0.304 24.168 ;
      RECT 0.000 22.192 0.304 22.952 ;
      RECT 0.000 20.976 0.304 21.736 ;
      RECT 0.000 19.760 0.304 20.520 ;
      RECT 0.000 18.544 0.304 19.304 ;
      RECT 0.000 17.328 0.304 18.088 ;
      RECT 0.000 16.112 0.304 16.872 ;
      RECT 0.000 14.896 0.304 15.656 ;
      RECT 0.000 0.304 0.304 14.440 ;
      RECT 0.000 134.040 5.043 136.192 ;
      RECT 7.355 134.040 7.763 136.192 ;
      RECT 10.067 134.040 278.464 136.192 ;
      RECT 0.304 0.304 278.160 134.040 ;
  END

END sram8t512x128

END LIBRARY
