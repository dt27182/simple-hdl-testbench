VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram6t4096x64
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 205.504 BY 358.720 ;
  SYMMETRY X Y R90 ;

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 195.168 0.000 195.320 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 195.168 0.000 195.320 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 195.168 0.000 195.320 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 195.168 0.000 195.320 0.152 ;
    END
  END CE1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 190.608 0.000 190.760 0.152 ;
    END
  END CSB1

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.048 0.000 186.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 186.048 0.000 186.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 186.048 0.000 186.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 186.048 0.000 186.200 0.152 ;
    END
  END OEB1

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 181.488 0.000 181.640 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 181.488 0.000 181.640 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 181.488 0.000 181.640 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 181.488 0.000 181.640 0.152 ;
    END
  END O1[3]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 181.184 0.000 181.336 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 181.184 0.000 181.336 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 181.184 0.000 181.336 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 181.184 0.000 181.336 0.152 ;
    END
  END O1[2]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 180.880 0.000 181.032 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 180.880 0.000 181.032 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 180.880 0.000 181.032 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 180.880 0.000 181.032 0.152 ;
    END
  END O1[1]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 180.576 0.000 180.728 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 180.576 0.000 180.728 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 180.576 0.000 180.728 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 180.576 0.000 180.728 0.152 ;
    END
  END O1[0]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.016 0.000 176.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 176.016 0.000 176.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 176.016 0.000 176.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 176.016 0.000 176.168 0.152 ;
    END
  END I1[0]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.712 0.000 175.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 175.712 0.000 175.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 175.712 0.000 175.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.712 0.000 175.864 0.152 ;
    END
  END I1[1]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.408 0.000 175.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 175.408 0.000 175.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 175.408 0.000 175.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.408 0.000 175.560 0.152 ;
    END
  END I1[2]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.104 0.000 175.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 175.104 0.000 175.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 175.104 0.000 175.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 175.104 0.000 175.256 0.152 ;
    END
  END I1[3]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.544 0.000 170.696 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 170.544 0.000 170.696 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 170.544 0.000 170.696 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 170.544 0.000 170.696 0.152 ;
    END
  END O1[7]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.240 0.000 170.392 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 170.240 0.000 170.392 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 170.240 0.000 170.392 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 170.240 0.000 170.392 0.152 ;
    END
  END O1[6]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 169.936 0.000 170.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 169.936 0.000 170.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 169.936 0.000 170.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 169.936 0.000 170.088 0.152 ;
    END
  END O1[5]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 169.632 0.000 169.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 169.632 0.000 169.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 169.632 0.000 169.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 169.632 0.000 169.784 0.152 ;
    END
  END O1[4]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.072 0.000 165.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 165.072 0.000 165.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 165.072 0.000 165.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 165.072 0.000 165.224 0.152 ;
    END
  END I1[4]

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.768 0.000 164.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 164.768 0.000 164.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 164.768 0.000 164.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 164.768 0.000 164.920 0.152 ;
    END
  END I1[5]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.464 0.000 164.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 164.464 0.000 164.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 164.464 0.000 164.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 164.464 0.000 164.616 0.152 ;
    END
  END I1[6]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.160 0.000 164.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 164.160 0.000 164.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 164.160 0.000 164.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 164.160 0.000 164.312 0.152 ;
    END
  END I1[7]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.600 0.000 159.752 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 159.600 0.000 159.752 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 159.600 0.000 159.752 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 159.600 0.000 159.752 0.152 ;
    END
  END O1[11]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.296 0.000 159.448 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 159.296 0.000 159.448 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 159.296 0.000 159.448 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 159.296 0.000 159.448 0.152 ;
    END
  END O1[10]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.992 0.000 159.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 158.992 0.000 159.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 158.992 0.000 159.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 158.992 0.000 159.144 0.152 ;
    END
  END O1[9]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.688 0.000 158.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 158.688 0.000 158.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 158.688 0.000 158.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 158.688 0.000 158.840 0.152 ;
    END
  END O1[8]

  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 154.128 0.000 154.280 0.152 ;
    END
  END I1[8]

  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.824 0.000 153.976 0.152 ;
    END
  END I1[9]

  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
  END I1[10]

  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
  END I1[11]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.656 0.000 148.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.656 0.000 148.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.656 0.000 148.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.656 0.000 148.808 0.152 ;
    END
  END O1[15]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.352 0.000 148.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.352 0.000 148.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.352 0.000 148.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.352 0.000 148.504 0.152 ;
    END
  END O1[14]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.048 0.000 148.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.048 0.000 148.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.048 0.000 148.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.048 0.000 148.200 0.152 ;
    END
  END O1[13]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.744 0.000 147.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 147.744 0.000 147.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 147.744 0.000 147.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 147.744 0.000 147.896 0.152 ;
    END
  END O1[12]

  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.184 0.000 143.336 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 143.184 0.000 143.336 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 143.184 0.000 143.336 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 143.184 0.000 143.336 0.152 ;
    END
  END I1[12]

  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.880 0.000 143.032 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 142.880 0.000 143.032 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 142.880 0.000 143.032 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 142.880 0.000 143.032 0.152 ;
    END
  END I1[13]

  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.576 0.000 142.728 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 142.576 0.000 142.728 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 142.576 0.000 142.728 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 142.576 0.000 142.728 0.152 ;
    END
  END I1[14]

  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.272 0.000 142.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 142.272 0.000 142.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 142.272 0.000 142.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 142.272 0.000 142.424 0.152 ;
    END
  END I1[15]

  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.712 0.000 137.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 137.712 0.000 137.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 137.712 0.000 137.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 137.712 0.000 137.864 0.152 ;
    END
  END O1[19]

  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.408 0.000 137.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 137.408 0.000 137.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 137.408 0.000 137.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 137.408 0.000 137.560 0.152 ;
    END
  END O1[18]

  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.104 0.000 137.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 137.104 0.000 137.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 137.104 0.000 137.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 137.104 0.000 137.256 0.152 ;
    END
  END O1[17]

  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.800 0.000 136.952 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 136.800 0.000 136.952 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 136.800 0.000 136.952 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 136.800 0.000 136.952 0.152 ;
    END
  END O1[16]

  PIN I1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.240 0.000 132.392 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.240 0.000 132.392 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.240 0.000 132.392 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 132.240 0.000 132.392 0.152 ;
    END
  END I1[16]

  PIN I1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.936 0.000 132.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.936 0.000 132.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.936 0.000 132.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.936 0.000 132.088 0.152 ;
    END
  END I1[17]

  PIN I1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.632 0.000 131.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.632 0.000 131.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.632 0.000 131.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.632 0.000 131.784 0.152 ;
    END
  END I1[18]

  PIN I1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.328 0.000 131.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.328 0.000 131.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.328 0.000 131.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.328 0.000 131.480 0.152 ;
    END
  END I1[19]

  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.768 0.000 126.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 126.768 0.000 126.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 126.768 0.000 126.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.768 0.000 126.920 0.152 ;
    END
  END O1[23]

  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.464 0.000 126.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 126.464 0.000 126.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 126.464 0.000 126.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.464 0.000 126.616 0.152 ;
    END
  END O1[22]

  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.160 0.000 126.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 126.160 0.000 126.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 126.160 0.000 126.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.160 0.000 126.312 0.152 ;
    END
  END O1[21]

  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.856 0.000 126.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 125.856 0.000 126.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 125.856 0.000 126.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.856 0.000 126.008 0.152 ;
    END
  END O1[20]

  PIN I1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.296 0.000 121.448 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 121.296 0.000 121.448 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 121.296 0.000 121.448 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.296 0.000 121.448 0.152 ;
    END
  END I1[20]

  PIN I1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.992 0.000 121.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.992 0.000 121.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.992 0.000 121.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.992 0.000 121.144 0.152 ;
    END
  END I1[21]

  PIN I1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.688 0.000 120.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.688 0.000 120.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.688 0.000 120.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.688 0.000 120.840 0.152 ;
    END
  END I1[22]

  PIN I1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.384 0.000 120.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.384 0.000 120.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.384 0.000 120.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.384 0.000 120.536 0.152 ;
    END
  END I1[23]

  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.824 0.000 115.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 115.824 0.000 115.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 115.824 0.000 115.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.824 0.000 115.976 0.152 ;
    END
  END O1[27]

  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.520 0.000 115.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 115.520 0.000 115.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 115.520 0.000 115.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.520 0.000 115.672 0.152 ;
    END
  END O1[26]

  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.216 0.000 115.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 115.216 0.000 115.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 115.216 0.000 115.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.216 0.000 115.368 0.152 ;
    END
  END O1[25]

  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.912 0.000 115.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 114.912 0.000 115.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 114.912 0.000 115.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.912 0.000 115.064 0.152 ;
    END
  END O1[24]

  PIN I1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.352 0.000 110.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.352 0.000 110.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.352 0.000 110.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.352 0.000 110.504 0.152 ;
    END
  END I1[24]

  PIN I1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
  END I1[25]

  PIN I1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.744 0.000 109.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.744 0.000 109.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.744 0.000 109.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.744 0.000 109.896 0.152 ;
    END
  END I1[26]

  PIN I1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.440 0.000 109.592 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.440 0.000 109.592 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.440 0.000 109.592 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.440 0.000 109.592 0.152 ;
    END
  END I1[27]

  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.880 0.000 105.032 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.880 0.000 105.032 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.880 0.000 105.032 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.880 0.000 105.032 0.152 ;
    END
  END O1[31]

  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.576 0.000 104.728 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.576 0.000 104.728 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.576 0.000 104.728 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.576 0.000 104.728 0.152 ;
    END
  END O1[30]

  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.272 0.000 104.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.272 0.000 104.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.272 0.000 104.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.272 0.000 104.424 0.152 ;
    END
  END O1[29]

  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.968 0.000 104.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.968 0.000 104.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.968 0.000 104.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.968 0.000 104.120 0.152 ;
    END
  END O1[28]

  PIN I1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.408 0.000 99.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.408 0.000 99.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.408 0.000 99.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.408 0.000 99.560 0.152 ;
    END
  END I1[28]

  PIN I1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.104 0.000 99.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.104 0.000 99.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.104 0.000 99.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.104 0.000 99.256 0.152 ;
    END
  END I1[29]

  PIN I1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.800 0.000 98.952 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.800 0.000 98.952 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.800 0.000 98.952 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.800 0.000 98.952 0.152 ;
    END
  END I1[30]

  PIN I1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.496 0.000 98.648 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.496 0.000 98.648 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.496 0.000 98.648 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.496 0.000 98.648 0.152 ;
    END
  END I1[31]

  PIN O1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.936 0.000 94.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.936 0.000 94.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.936 0.000 94.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.936 0.000 94.088 0.152 ;
    END
  END O1[35]

  PIN O1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.632 0.000 93.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.632 0.000 93.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.632 0.000 93.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.632 0.000 93.784 0.152 ;
    END
  END O1[34]

  PIN O1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.328 0.000 93.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.328 0.000 93.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.328 0.000 93.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.328 0.000 93.480 0.152 ;
    END
  END O1[33]

  PIN O1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
  END O1[32]

  PIN I1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.464 0.000 88.616 0.152 ;
    END
  END I1[32]

  PIN I1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.160 0.000 88.312 0.152 ;
    END
  END I1[33]

  PIN I1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.856 0.000 88.008 0.152 ;
    END
  END I1[34]

  PIN I1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.552 0.000 87.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.552 0.000 87.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.552 0.000 87.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.552 0.000 87.704 0.152 ;
    END
  END I1[35]

  PIN O1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.992 0.000 83.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.992 0.000 83.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.992 0.000 83.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.992 0.000 83.144 0.152 ;
    END
  END O1[39]

  PIN O1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.688 0.000 82.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.688 0.000 82.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.688 0.000 82.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.688 0.000 82.840 0.152 ;
    END
  END O1[38]

  PIN O1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
  END O1[37]

  PIN O1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.080 0.000 82.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.080 0.000 82.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.080 0.000 82.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.080 0.000 82.232 0.152 ;
    END
  END O1[36]

  PIN I1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.520 0.000 77.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.520 0.000 77.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.520 0.000 77.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.520 0.000 77.672 0.152 ;
    END
  END I1[36]

  PIN I1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.216 0.000 77.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 77.216 0.000 77.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 77.216 0.000 77.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 77.216 0.000 77.368 0.152 ;
    END
  END I1[37]

  PIN I1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.912 0.000 77.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.912 0.000 77.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.912 0.000 77.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.912 0.000 77.064 0.152 ;
    END
  END I1[38]

  PIN I1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.608 0.000 76.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.608 0.000 76.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.608 0.000 76.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.608 0.000 76.760 0.152 ;
    END
  END I1[39]

  PIN O1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.048 0.000 72.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.048 0.000 72.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.048 0.000 72.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.048 0.000 72.200 0.152 ;
    END
  END O1[43]

  PIN O1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
  END O1[42]

  PIN O1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.440 0.000 71.592 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.440 0.000 71.592 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.440 0.000 71.592 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.440 0.000 71.592 0.152 ;
    END
  END O1[41]

  PIN O1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.136 0.000 71.288 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.136 0.000 71.288 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.136 0.000 71.288 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.136 0.000 71.288 0.152 ;
    END
  END O1[40]

  PIN I1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.576 0.000 66.728 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.576 0.000 66.728 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.576 0.000 66.728 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.576 0.000 66.728 0.152 ;
    END
  END I1[40]

  PIN I1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.272 0.000 66.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.272 0.000 66.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.272 0.000 66.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.272 0.000 66.424 0.152 ;
    END
  END I1[41]

  PIN I1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.968 0.000 66.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.968 0.000 66.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.968 0.000 66.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.968 0.000 66.120 0.152 ;
    END
  END I1[42]

  PIN I1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.664 0.000 65.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.664 0.000 65.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.664 0.000 65.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.664 0.000 65.816 0.152 ;
    END
  END I1[43]

  PIN O1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.104 0.000 61.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.104 0.000 61.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.104 0.000 61.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.104 0.000 61.256 0.152 ;
    END
  END O1[47]

  PIN O1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.800 0.000 60.952 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.800 0.000 60.952 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.800 0.000 60.952 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.800 0.000 60.952 0.152 ;
    END
  END O1[46]

  PIN O1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.496 0.000 60.648 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.496 0.000 60.648 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.496 0.000 60.648 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.496 0.000 60.648 0.152 ;
    END
  END O1[45]

  PIN O1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.192 0.000 60.344 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.192 0.000 60.344 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.192 0.000 60.344 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.192 0.000 60.344 0.152 ;
    END
  END O1[44]

  PIN I1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.632 0.000 55.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.632 0.000 55.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.632 0.000 55.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.632 0.000 55.784 0.152 ;
    END
  END I1[44]

  PIN I1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.328 0.000 55.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.328 0.000 55.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.328 0.000 55.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.328 0.000 55.480 0.152 ;
    END
  END I1[45]

  PIN I1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.024 0.000 55.176 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.024 0.000 55.176 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.024 0.000 55.176 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.024 0.000 55.176 0.152 ;
    END
  END I1[46]

  PIN I1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.720 0.000 54.872 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.720 0.000 54.872 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.720 0.000 54.872 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.720 0.000 54.872 0.152 ;
    END
  END I1[47]

  PIN O1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
  END O1[51]

  PIN O1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
  END O1[50]

  PIN O1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.552 0.000 49.704 0.152 ;
    END
  END O1[49]

  PIN O1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
  END O1[48]

  PIN I1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
  END I1[48]

  PIN I1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.384 0.000 44.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.384 0.000 44.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.384 0.000 44.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.384 0.000 44.536 0.152 ;
    END
  END I1[49]

  PIN I1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
  END I1[50]

  PIN I1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.776 0.000 43.928 0.152 ;
    END
  END I1[51]

  PIN O1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
  END O1[55]

  PIN O1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
  END O1[54]

  PIN O1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
  END O1[53]

  PIN O1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
  END O1[52]

  PIN I1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.744 0.000 33.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.744 0.000 33.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.744 0.000 33.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.744 0.000 33.896 0.152 ;
    END
  END I1[52]

  PIN I1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.440 0.000 33.592 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.440 0.000 33.592 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.440 0.000 33.592 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.440 0.000 33.592 0.152 ;
    END
  END I1[53]

  PIN I1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.136 0.000 33.288 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.136 0.000 33.288 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.136 0.000 33.288 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.136 0.000 33.288 0.152 ;
    END
  END I1[54]

  PIN I1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.832 0.000 32.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.832 0.000 32.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.832 0.000 32.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.832 0.000 32.984 0.152 ;
    END
  END I1[55]

  PIN O1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.272 0.000 28.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.272 0.000 28.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.272 0.000 28.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.272 0.000 28.424 0.152 ;
    END
  END O1[59]

  PIN O1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
  END O1[58]

  PIN O1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.664 0.000 27.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.664 0.000 27.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.664 0.000 27.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.664 0.000 27.816 0.152 ;
    END
  END O1[57]

  PIN O1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.360 0.000 27.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.360 0.000 27.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.360 0.000 27.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.360 0.000 27.512 0.152 ;
    END
  END O1[56]

  PIN I1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.800 0.000 22.952 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.800 0.000 22.952 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.800 0.000 22.952 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.800 0.000 22.952 0.152 ;
    END
  END I1[56]

  PIN I1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.496 0.000 22.648 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.496 0.000 22.648 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.496 0.000 22.648 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.496 0.000 22.648 0.152 ;
    END
  END I1[57]

  PIN I1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.192 0.000 22.344 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.192 0.000 22.344 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.192 0.000 22.344 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.192 0.000 22.344 0.152 ;
    END
  END I1[58]

  PIN I1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.888 0.000 22.040 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.888 0.000 22.040 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.888 0.000 22.040 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.888 0.000 22.040 0.152 ;
    END
  END I1[59]

  PIN O1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.328 0.000 17.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.328 0.000 17.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.328 0.000 17.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.328 0.000 17.480 0.152 ;
    END
  END O1[63]

  PIN O1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.024 0.000 17.176 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.024 0.000 17.176 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.024 0.000 17.176 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.024 0.000 17.176 0.152 ;
    END
  END O1[62]

  PIN O1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.720 0.000 16.872 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.720 0.000 16.872 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.720 0.000 16.872 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.720 0.000 16.872 0.152 ;
    END
  END O1[61]

  PIN O1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.416 0.000 16.568 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 16.416 0.000 16.568 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 16.416 0.000 16.568 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 16.416 0.000 16.568 0.152 ;
    END
  END O1[60]

  PIN I1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.856 0.000 12.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.856 0.000 12.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.856 0.000 12.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.856 0.000 12.008 0.152 ;
    END
  END I1[60]

  PIN I1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.552 0.000 11.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.552 0.000 11.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.552 0.000 11.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.552 0.000 11.704 0.152 ;
    END
  END I1[61]

  PIN I1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.248 0.000 11.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 11.248 0.000 11.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 11.248 0.000 11.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 11.248 0.000 11.400 0.152 ;
    END
  END I1[62]

  PIN I1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.944 0.000 11.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.944 0.000 11.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.944 0.000 11.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.944 0.000 11.096 0.152 ;
    END
  END I1[63]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 313.880 205.504 314.032 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 313.880 205.504 314.032 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 313.880 205.504 314.032 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 313.880 205.504 314.032 ;
    END
  END A1[0]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 310.232 205.504 310.384 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 310.232 205.504 310.384 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 310.232 205.504 310.384 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 310.232 205.504 310.384 ;
    END
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 306.584 205.504 306.736 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 306.584 205.504 306.736 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 306.584 205.504 306.736 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 306.584 205.504 306.736 ;
    END
  END A1[2]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 302.936 205.504 303.088 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 302.936 205.504 303.088 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 302.936 205.504 303.088 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 302.936 205.504 303.088 ;
    END
  END A1[3]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 299.288 205.504 299.440 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 299.288 205.504 299.440 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 299.288 205.504 299.440 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 299.288 205.504 299.440 ;
    END
  END A1[4]

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 295.640 205.504 295.792 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 295.640 205.504 295.792 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 295.640 205.504 295.792 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 295.640 205.504 295.792 ;
    END
  END A1[5]

  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 291.992 205.504 292.144 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 291.992 205.504 292.144 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 291.992 205.504 292.144 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 291.992 205.504 292.144 ;
    END
  END A1[6]

  PIN A1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 288.344 205.504 288.496 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 288.344 205.504 288.496 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 288.344 205.504 288.496 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 288.344 205.504 288.496 ;
    END
  END A1[7]

  PIN A1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 284.696 205.504 284.848 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 284.696 205.504 284.848 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 284.696 205.504 284.848 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 284.696 205.504 284.848 ;
    END
  END A1[8]

  PIN A1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 281.048 205.504 281.200 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 281.048 205.504 281.200 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 281.048 205.504 281.200 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 281.048 205.504 281.200 ;
    END
  END A1[9]

  PIN A1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 277.400 205.504 277.552 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 277.400 205.504 277.552 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 277.400 205.504 277.552 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 277.400 205.504 277.552 ;
    END
  END A1[10]

  PIN A1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 273.752 205.504 273.904 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 273.752 205.504 273.904 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 273.752 205.504 273.904 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 273.752 205.504 273.904 ;
    END
  END A1[11]

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 89.680 205.504 89.832 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 89.680 205.504 89.832 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 89.680 205.504 89.832 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 89.680 205.504 89.832 ;
    END
  END WEB1

  PIN WBM1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 88.464 205.504 88.616 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 88.464 205.504 88.616 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 88.464 205.504 88.616 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 88.464 205.504 88.616 ;
    END
  END WBM1[0]

  PIN WBM1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 87.248 205.504 87.400 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 87.248 205.504 87.400 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 87.248 205.504 87.400 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 87.248 205.504 87.400 ;
    END
  END WBM1[1]

  PIN WBM1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 86.032 205.504 86.184 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 86.032 205.504 86.184 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 86.032 205.504 86.184 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 86.032 205.504 86.184 ;
    END
  END WBM1[2]

  PIN WBM1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 84.816 205.504 84.968 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 84.816 205.504 84.968 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 84.816 205.504 84.968 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 84.816 205.504 84.968 ;
    END
  END WBM1[3]

  PIN WBM1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 83.600 205.504 83.752 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 83.600 205.504 83.752 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 83.600 205.504 83.752 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 83.600 205.504 83.752 ;
    END
  END WBM1[4]

  PIN WBM1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 82.384 205.504 82.536 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 82.384 205.504 82.536 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 82.384 205.504 82.536 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 82.384 205.504 82.536 ;
    END
  END WBM1[5]

  PIN WBM1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 81.168 205.504 81.320 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 81.168 205.504 81.320 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 81.168 205.504 81.320 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 81.168 205.504 81.320 ;
    END
  END WBM1[6]

  PIN WBM1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.352 79.952 205.504 80.104 ;
    END
    PORT
      LAYER M3 ;
        RECT 205.352 79.952 205.504 80.104 ;
    END
    PORT
      LAYER M4 ;
        RECT 205.352 79.952 205.504 80.104 ;
    END
    PORT
      LAYER M5 ;
        RECT 205.352 79.952 205.504 80.104 ;
    END
  END WBM1[7]

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 5.195 356.720 7.195 358.720 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.195 356.720 7.195 358.720 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.195 356.720 7.195 358.720 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M2 ;
        RECT 7.915 356.720 9.915 358.720 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.915 356.720 9.915 358.720 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.915 356.720 9.915 358.720 ;
    END
  END VSS

  OBS
    LAYER M2 ;
      RECT 195.472 0.000 205.504 0.304 ;
      RECT 190.912 0.000 195.016 0.304 ;
      RECT 186.352 0.000 190.456 0.304 ;
      RECT 181.792 0.000 185.896 0.304 ;
      RECT 176.320 0.000 180.424 0.304 ;
      RECT 170.848 0.000 174.952 0.304 ;
      RECT 165.376 0.000 169.480 0.304 ;
      RECT 159.904 0.000 164.008 0.304 ;
      RECT 154.432 0.000 158.536 0.304 ;
      RECT 148.960 0.000 153.064 0.304 ;
      RECT 143.488 0.000 147.592 0.304 ;
      RECT 138.016 0.000 142.120 0.304 ;
      RECT 132.544 0.000 136.648 0.304 ;
      RECT 127.072 0.000 131.176 0.304 ;
      RECT 121.600 0.000 125.704 0.304 ;
      RECT 116.128 0.000 120.232 0.304 ;
      RECT 110.656 0.000 114.760 0.304 ;
      RECT 105.184 0.000 109.288 0.304 ;
      RECT 99.712 0.000 103.816 0.304 ;
      RECT 94.240 0.000 98.344 0.304 ;
      RECT 88.768 0.000 92.872 0.304 ;
      RECT 83.296 0.000 87.400 0.304 ;
      RECT 77.824 0.000 81.928 0.304 ;
      RECT 72.352 0.000 76.456 0.304 ;
      RECT 66.880 0.000 70.984 0.304 ;
      RECT 61.408 0.000 65.512 0.304 ;
      RECT 55.936 0.000 60.040 0.304 ;
      RECT 50.464 0.000 54.568 0.304 ;
      RECT 44.992 0.000 49.096 0.304 ;
      RECT 39.520 0.000 43.624 0.304 ;
      RECT 34.048 0.000 38.152 0.304 ;
      RECT 28.576 0.000 32.680 0.304 ;
      RECT 23.104 0.000 27.208 0.304 ;
      RECT 17.632 0.000 21.736 0.304 ;
      RECT 12.160 0.000 16.264 0.304 ;
      RECT 0.000 0.000 10.792 0.304 ;
      RECT 205.200 314.184 205.504 356.568 ;
      RECT 205.200 310.536 205.504 313.728 ;
      RECT 205.200 306.888 205.504 310.080 ;
      RECT 205.200 303.240 205.504 306.432 ;
      RECT 205.200 299.592 205.504 302.784 ;
      RECT 205.200 295.944 205.504 299.136 ;
      RECT 205.200 292.296 205.504 295.488 ;
      RECT 205.200 288.648 205.504 291.840 ;
      RECT 205.200 285.000 205.504 288.192 ;
      RECT 205.200 281.352 205.504 284.544 ;
      RECT 205.200 277.704 205.504 280.896 ;
      RECT 205.200 274.056 205.504 277.248 ;
      RECT 205.200 89.984 205.504 273.600 ;
      RECT 205.200 88.768 205.504 89.528 ;
      RECT 205.200 87.552 205.504 88.312 ;
      RECT 205.200 86.336 205.504 87.096 ;
      RECT 205.200 85.120 205.504 85.880 ;
      RECT 205.200 83.904 205.504 84.664 ;
      RECT 205.200 82.688 205.504 83.448 ;
      RECT 205.200 81.472 205.504 82.232 ;
      RECT 205.200 80.256 205.504 81.016 ;
      RECT 205.200 0.304 205.504 79.800 ;
      RECT 0.000 356.568 5.043 358.720 ;
      RECT 7.355 356.568 7.763 358.720 ;
      RECT 10.067 356.568 205.504 358.720 ;
      RECT 0.000 0.304 205.200 356.568 ;
    LAYER M3 ;
      RECT 195.472 0.000 205.504 0.304 ;
      RECT 190.912 0.000 195.016 0.304 ;
      RECT 186.352 0.000 190.456 0.304 ;
      RECT 181.792 0.000 185.896 0.304 ;
      RECT 176.320 0.000 180.424 0.304 ;
      RECT 170.848 0.000 174.952 0.304 ;
      RECT 165.376 0.000 169.480 0.304 ;
      RECT 159.904 0.000 164.008 0.304 ;
      RECT 154.432 0.000 158.536 0.304 ;
      RECT 148.960 0.000 153.064 0.304 ;
      RECT 143.488 0.000 147.592 0.304 ;
      RECT 138.016 0.000 142.120 0.304 ;
      RECT 132.544 0.000 136.648 0.304 ;
      RECT 127.072 0.000 131.176 0.304 ;
      RECT 121.600 0.000 125.704 0.304 ;
      RECT 116.128 0.000 120.232 0.304 ;
      RECT 110.656 0.000 114.760 0.304 ;
      RECT 105.184 0.000 109.288 0.304 ;
      RECT 99.712 0.000 103.816 0.304 ;
      RECT 94.240 0.000 98.344 0.304 ;
      RECT 88.768 0.000 92.872 0.304 ;
      RECT 83.296 0.000 87.400 0.304 ;
      RECT 77.824 0.000 81.928 0.304 ;
      RECT 72.352 0.000 76.456 0.304 ;
      RECT 66.880 0.000 70.984 0.304 ;
      RECT 61.408 0.000 65.512 0.304 ;
      RECT 55.936 0.000 60.040 0.304 ;
      RECT 50.464 0.000 54.568 0.304 ;
      RECT 44.992 0.000 49.096 0.304 ;
      RECT 39.520 0.000 43.624 0.304 ;
      RECT 34.048 0.000 38.152 0.304 ;
      RECT 28.576 0.000 32.680 0.304 ;
      RECT 23.104 0.000 27.208 0.304 ;
      RECT 17.632 0.000 21.736 0.304 ;
      RECT 12.160 0.000 16.264 0.304 ;
      RECT 0.000 0.000 10.792 0.304 ;
      RECT 205.200 314.184 205.504 356.568 ;
      RECT 205.200 310.536 205.504 313.728 ;
      RECT 205.200 306.888 205.504 310.080 ;
      RECT 205.200 303.240 205.504 306.432 ;
      RECT 205.200 299.592 205.504 302.784 ;
      RECT 205.200 295.944 205.504 299.136 ;
      RECT 205.200 292.296 205.504 295.488 ;
      RECT 205.200 288.648 205.504 291.840 ;
      RECT 205.200 285.000 205.504 288.192 ;
      RECT 205.200 281.352 205.504 284.544 ;
      RECT 205.200 277.704 205.504 280.896 ;
      RECT 205.200 274.056 205.504 277.248 ;
      RECT 205.200 89.984 205.504 273.600 ;
      RECT 205.200 88.768 205.504 89.528 ;
      RECT 205.200 87.552 205.504 88.312 ;
      RECT 205.200 86.336 205.504 87.096 ;
      RECT 205.200 85.120 205.504 85.880 ;
      RECT 205.200 83.904 205.504 84.664 ;
      RECT 205.200 82.688 205.504 83.448 ;
      RECT 205.200 81.472 205.504 82.232 ;
      RECT 205.200 80.256 205.504 81.016 ;
      RECT 205.200 0.304 205.504 79.800 ;
      RECT 0.000 356.568 5.043 358.720 ;
      RECT 7.355 356.568 7.763 358.720 ;
      RECT 10.067 356.568 205.504 358.720 ;
      RECT 0.000 0.304 205.200 356.568 ;
    LAYER M4 ;
      RECT 195.472 0.000 205.504 0.304 ;
      RECT 190.912 0.000 195.016 0.304 ;
      RECT 186.352 0.000 190.456 0.304 ;
      RECT 181.792 0.000 185.896 0.304 ;
      RECT 176.320 0.000 180.424 0.304 ;
      RECT 170.848 0.000 174.952 0.304 ;
      RECT 165.376 0.000 169.480 0.304 ;
      RECT 159.904 0.000 164.008 0.304 ;
      RECT 154.432 0.000 158.536 0.304 ;
      RECT 148.960 0.000 153.064 0.304 ;
      RECT 143.488 0.000 147.592 0.304 ;
      RECT 138.016 0.000 142.120 0.304 ;
      RECT 132.544 0.000 136.648 0.304 ;
      RECT 127.072 0.000 131.176 0.304 ;
      RECT 121.600 0.000 125.704 0.304 ;
      RECT 116.128 0.000 120.232 0.304 ;
      RECT 110.656 0.000 114.760 0.304 ;
      RECT 105.184 0.000 109.288 0.304 ;
      RECT 99.712 0.000 103.816 0.304 ;
      RECT 94.240 0.000 98.344 0.304 ;
      RECT 88.768 0.000 92.872 0.304 ;
      RECT 83.296 0.000 87.400 0.304 ;
      RECT 77.824 0.000 81.928 0.304 ;
      RECT 72.352 0.000 76.456 0.304 ;
      RECT 66.880 0.000 70.984 0.304 ;
      RECT 61.408 0.000 65.512 0.304 ;
      RECT 55.936 0.000 60.040 0.304 ;
      RECT 50.464 0.000 54.568 0.304 ;
      RECT 44.992 0.000 49.096 0.304 ;
      RECT 39.520 0.000 43.624 0.304 ;
      RECT 34.048 0.000 38.152 0.304 ;
      RECT 28.576 0.000 32.680 0.304 ;
      RECT 23.104 0.000 27.208 0.304 ;
      RECT 17.632 0.000 21.736 0.304 ;
      RECT 12.160 0.000 16.264 0.304 ;
      RECT 0.000 0.000 10.792 0.304 ;
      RECT 205.200 314.184 205.504 356.568 ;
      RECT 205.200 310.536 205.504 313.728 ;
      RECT 205.200 306.888 205.504 310.080 ;
      RECT 205.200 303.240 205.504 306.432 ;
      RECT 205.200 299.592 205.504 302.784 ;
      RECT 205.200 295.944 205.504 299.136 ;
      RECT 205.200 292.296 205.504 295.488 ;
      RECT 205.200 288.648 205.504 291.840 ;
      RECT 205.200 285.000 205.504 288.192 ;
      RECT 205.200 281.352 205.504 284.544 ;
      RECT 205.200 277.704 205.504 280.896 ;
      RECT 205.200 274.056 205.504 277.248 ;
      RECT 205.200 89.984 205.504 273.600 ;
      RECT 205.200 88.768 205.504 89.528 ;
      RECT 205.200 87.552 205.504 88.312 ;
      RECT 205.200 86.336 205.504 87.096 ;
      RECT 205.200 85.120 205.504 85.880 ;
      RECT 205.200 83.904 205.504 84.664 ;
      RECT 205.200 82.688 205.504 83.448 ;
      RECT 205.200 81.472 205.504 82.232 ;
      RECT 205.200 80.256 205.504 81.016 ;
      RECT 205.200 0.304 205.504 79.800 ;
      RECT 0.000 356.568 5.043 358.720 ;
      RECT 7.355 356.568 7.763 358.720 ;
      RECT 10.067 356.568 205.504 358.720 ;
      RECT 0.000 0.304 205.200 356.568 ;
    LAYER M5 ;
      RECT 195.472 0.000 205.504 0.304 ;
      RECT 190.912 0.000 195.016 0.304 ;
      RECT 186.352 0.000 190.456 0.304 ;
      RECT 181.792 0.000 185.896 0.304 ;
      RECT 176.320 0.000 180.424 0.304 ;
      RECT 170.848 0.000 174.952 0.304 ;
      RECT 165.376 0.000 169.480 0.304 ;
      RECT 159.904 0.000 164.008 0.304 ;
      RECT 154.432 0.000 158.536 0.304 ;
      RECT 148.960 0.000 153.064 0.304 ;
      RECT 143.488 0.000 147.592 0.304 ;
      RECT 138.016 0.000 142.120 0.304 ;
      RECT 132.544 0.000 136.648 0.304 ;
      RECT 127.072 0.000 131.176 0.304 ;
      RECT 121.600 0.000 125.704 0.304 ;
      RECT 116.128 0.000 120.232 0.304 ;
      RECT 110.656 0.000 114.760 0.304 ;
      RECT 105.184 0.000 109.288 0.304 ;
      RECT 99.712 0.000 103.816 0.304 ;
      RECT 94.240 0.000 98.344 0.304 ;
      RECT 88.768 0.000 92.872 0.304 ;
      RECT 83.296 0.000 87.400 0.304 ;
      RECT 77.824 0.000 81.928 0.304 ;
      RECT 72.352 0.000 76.456 0.304 ;
      RECT 66.880 0.000 70.984 0.304 ;
      RECT 61.408 0.000 65.512 0.304 ;
      RECT 55.936 0.000 60.040 0.304 ;
      RECT 50.464 0.000 54.568 0.304 ;
      RECT 44.992 0.000 49.096 0.304 ;
      RECT 39.520 0.000 43.624 0.304 ;
      RECT 34.048 0.000 38.152 0.304 ;
      RECT 28.576 0.000 32.680 0.304 ;
      RECT 23.104 0.000 27.208 0.304 ;
      RECT 17.632 0.000 21.736 0.304 ;
      RECT 12.160 0.000 16.264 0.304 ;
      RECT 0.000 0.000 10.792 0.304 ;
      RECT 205.200 314.184 205.504 356.568 ;
      RECT 205.200 310.536 205.504 313.728 ;
      RECT 205.200 306.888 205.504 310.080 ;
      RECT 205.200 303.240 205.504 306.432 ;
      RECT 205.200 299.592 205.504 302.784 ;
      RECT 205.200 295.944 205.504 299.136 ;
      RECT 205.200 292.296 205.504 295.488 ;
      RECT 205.200 288.648 205.504 291.840 ;
      RECT 205.200 285.000 205.504 288.192 ;
      RECT 205.200 281.352 205.504 284.544 ;
      RECT 205.200 277.704 205.504 280.896 ;
      RECT 205.200 274.056 205.504 277.248 ;
      RECT 205.200 89.984 205.504 273.600 ;
      RECT 205.200 88.768 205.504 89.528 ;
      RECT 205.200 87.552 205.504 88.312 ;
      RECT 205.200 86.336 205.504 87.096 ;
      RECT 205.200 85.120 205.504 85.880 ;
      RECT 205.200 83.904 205.504 84.664 ;
      RECT 205.200 82.688 205.504 83.448 ;
      RECT 205.200 81.472 205.504 82.232 ;
      RECT 205.200 80.256 205.504 81.016 ;
      RECT 205.200 0.304 205.504 79.800 ;
      RECT 0.000 356.568 5.043 358.720 ;
      RECT 7.355 356.568 7.763 358.720 ;
      RECT 10.067 356.568 205.504 358.720 ;
      RECT 0.000 0.304 205.200 356.568 ;
  END

END sram6t4096x64

END LIBRARY
