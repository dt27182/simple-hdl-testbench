VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram8t256x72
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 161.728 BY 74.176 ;
  SYMMETRY X Y R90 ;

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.472 0.000 157.624 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 157.472 0.000 157.624 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 157.472 0.000 157.624 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 157.472 0.000 157.624 0.152 ;
    END
  END CE1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.736 0.000 154.888 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.736 0.000 154.888 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.736 0.000 154.888 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 154.736 0.000 154.888 0.152 ;
    END
  END CSB1

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.000 0.000 152.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 152.000 0.000 152.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 152.000 0.000 152.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 152.000 0.000 152.152 0.152 ;
    END
  END OEB1

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.264 0.000 149.416 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 149.264 0.000 149.416 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 149.264 0.000 149.416 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 149.264 0.000 149.416 0.152 ;
    END
  END O1[3]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.960 0.000 149.112 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.960 0.000 149.112 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.960 0.000 149.112 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.960 0.000 149.112 0.152 ;
    END
  END O1[2]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.656 0.000 148.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.656 0.000 148.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.656 0.000 148.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.656 0.000 148.808 0.152 ;
    END
  END O1[1]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.352 0.000 148.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.352 0.000 148.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.352 0.000 148.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.352 0.000 148.504 0.152 ;
    END
  END O1[0]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.616 0.000 145.768 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 145.616 0.000 145.768 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 145.616 0.000 145.768 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.616 0.000 145.768 0.152 ;
    END
  END O1[7]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.312 0.000 145.464 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 145.312 0.000 145.464 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 145.312 0.000 145.464 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.312 0.000 145.464 0.152 ;
    END
  END O1[6]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.008 0.000 145.160 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 145.008 0.000 145.160 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 145.008 0.000 145.160 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.008 0.000 145.160 0.152 ;
    END
  END O1[5]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.704 0.000 144.856 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 144.704 0.000 144.856 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 144.704 0.000 144.856 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 144.704 0.000 144.856 0.152 ;
    END
  END O1[4]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.968 0.000 142.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 141.968 0.000 142.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.968 0.000 142.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.968 0.000 142.120 0.152 ;
    END
  END O1[11]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.664 0.000 141.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 141.664 0.000 141.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.664 0.000 141.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.664 0.000 141.816 0.152 ;
    END
  END O1[10]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.360 0.000 141.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 141.360 0.000 141.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.360 0.000 141.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.360 0.000 141.512 0.152 ;
    END
  END O1[9]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.056 0.000 141.208 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 141.056 0.000 141.208 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.056 0.000 141.208 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.056 0.000 141.208 0.152 ;
    END
  END O1[8]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.320 0.000 138.472 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 138.320 0.000 138.472 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 138.320 0.000 138.472 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 138.320 0.000 138.472 0.152 ;
    END
  END O1[15]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.016 0.000 138.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 138.016 0.000 138.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 138.016 0.000 138.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 138.016 0.000 138.168 0.152 ;
    END
  END O1[14]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.712 0.000 137.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 137.712 0.000 137.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 137.712 0.000 137.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 137.712 0.000 137.864 0.152 ;
    END
  END O1[13]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.408 0.000 137.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 137.408 0.000 137.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 137.408 0.000 137.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 137.408 0.000 137.560 0.152 ;
    END
  END O1[12]

  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.672 0.000 134.824 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 134.672 0.000 134.824 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 134.672 0.000 134.824 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.672 0.000 134.824 0.152 ;
    END
  END O1[19]

  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.368 0.000 134.520 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 134.368 0.000 134.520 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 134.368 0.000 134.520 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.368 0.000 134.520 0.152 ;
    END
  END O1[18]

  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.064 0.000 134.216 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 134.064 0.000 134.216 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 134.064 0.000 134.216 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.064 0.000 134.216 0.152 ;
    END
  END O1[17]

  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.760 0.000 133.912 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 133.760 0.000 133.912 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 133.760 0.000 133.912 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 133.760 0.000 133.912 0.152 ;
    END
  END O1[16]

  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.024 0.000 131.176 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.024 0.000 131.176 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.024 0.000 131.176 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.024 0.000 131.176 0.152 ;
    END
  END O1[23]

  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.720 0.000 130.872 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 130.720 0.000 130.872 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 130.720 0.000 130.872 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.720 0.000 130.872 0.152 ;
    END
  END O1[22]

  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.416 0.000 130.568 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 130.416 0.000 130.568 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 130.416 0.000 130.568 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.416 0.000 130.568 0.152 ;
    END
  END O1[21]

  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.112 0.000 130.264 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 130.112 0.000 130.264 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 130.112 0.000 130.264 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.112 0.000 130.264 0.152 ;
    END
  END O1[20]

  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.376 0.000 127.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 127.376 0.000 127.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 127.376 0.000 127.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.376 0.000 127.528 0.152 ;
    END
  END O1[27]

  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.072 0.000 127.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 127.072 0.000 127.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 127.072 0.000 127.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.072 0.000 127.224 0.152 ;
    END
  END O1[26]

  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.768 0.000 126.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 126.768 0.000 126.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 126.768 0.000 126.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.768 0.000 126.920 0.152 ;
    END
  END O1[25]

  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 126.464 0.000 126.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 126.464 0.000 126.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 126.464 0.000 126.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 126.464 0.000 126.616 0.152 ;
    END
  END O1[24]

  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.728 0.000 123.880 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 123.728 0.000 123.880 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 123.728 0.000 123.880 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.728 0.000 123.880 0.152 ;
    END
  END O1[31]

  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.424 0.000 123.576 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 123.424 0.000 123.576 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 123.424 0.000 123.576 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.424 0.000 123.576 0.152 ;
    END
  END O1[30]

  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.120 0.000 123.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 123.120 0.000 123.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 123.120 0.000 123.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.120 0.000 123.272 0.152 ;
    END
  END O1[29]

  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.816 0.000 122.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 122.816 0.000 122.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 122.816 0.000 122.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.816 0.000 122.968 0.152 ;
    END
  END O1[28]

  PIN O1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.080 0.000 120.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.080 0.000 120.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.080 0.000 120.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.080 0.000 120.232 0.152 ;
    END
  END O1[35]

  PIN O1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.776 0.000 119.928 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 119.776 0.000 119.928 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 119.776 0.000 119.928 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.776 0.000 119.928 0.152 ;
    END
  END O1[34]

  PIN O1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.472 0.000 119.624 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 119.472 0.000 119.624 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 119.472 0.000 119.624 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.472 0.000 119.624 0.152 ;
    END
  END O1[33]

  PIN O1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.168 0.000 119.320 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 119.168 0.000 119.320 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 119.168 0.000 119.320 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.168 0.000 119.320 0.152 ;
    END
  END O1[32]

  PIN O1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.432 0.000 116.584 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 116.432 0.000 116.584 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 116.432 0.000 116.584 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.432 0.000 116.584 0.152 ;
    END
  END O1[39]

  PIN O1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.128 0.000 116.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 116.128 0.000 116.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 116.128 0.000 116.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.128 0.000 116.280 0.152 ;
    END
  END O1[38]

  PIN O1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.824 0.000 115.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 115.824 0.000 115.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 115.824 0.000 115.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.824 0.000 115.976 0.152 ;
    END
  END O1[37]

  PIN O1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.520 0.000 115.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 115.520 0.000 115.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 115.520 0.000 115.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.520 0.000 115.672 0.152 ;
    END
  END O1[36]

  PIN O1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.784 0.000 112.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 112.784 0.000 112.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.784 0.000 112.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.784 0.000 112.936 0.152 ;
    END
  END O1[43]

  PIN O1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.480 0.000 112.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 112.480 0.000 112.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.480 0.000 112.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.480 0.000 112.632 0.152 ;
    END
  END O1[42]

  PIN O1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.176 0.000 112.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 112.176 0.000 112.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.176 0.000 112.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.176 0.000 112.328 0.152 ;
    END
  END O1[41]

  PIN O1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.872 0.000 112.024 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 111.872 0.000 112.024 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 111.872 0.000 112.024 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 111.872 0.000 112.024 0.152 ;
    END
  END O1[40]

  PIN O1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.136 0.000 109.288 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 109.136 0.000 109.288 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 109.136 0.000 109.288 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 109.136 0.000 109.288 0.152 ;
    END
  END O1[47]

  PIN O1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.832 0.000 108.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.832 0.000 108.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.832 0.000 108.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.832 0.000 108.984 0.152 ;
    END
  END O1[46]

  PIN O1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.528 0.000 108.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.528 0.000 108.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.528 0.000 108.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.528 0.000 108.680 0.152 ;
    END
  END O1[45]

  PIN O1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.224 0.000 108.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.224 0.000 108.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.224 0.000 108.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.224 0.000 108.376 0.152 ;
    END
  END O1[44]

  PIN O1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.488 0.000 105.640 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.488 0.000 105.640 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.488 0.000 105.640 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.488 0.000 105.640 0.152 ;
    END
  END O1[51]

  PIN O1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.184 0.000 105.336 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.184 0.000 105.336 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.184 0.000 105.336 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.184 0.000 105.336 0.152 ;
    END
  END O1[50]

  PIN O1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.880 0.000 105.032 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.880 0.000 105.032 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.880 0.000 105.032 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.880 0.000 105.032 0.152 ;
    END
  END O1[49]

  PIN O1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.576 0.000 104.728 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.576 0.000 104.728 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.576 0.000 104.728 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.576 0.000 104.728 0.152 ;
    END
  END O1[48]

  PIN O1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.840 0.000 101.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.840 0.000 101.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.840 0.000 101.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.840 0.000 101.992 0.152 ;
    END
  END O1[55]

  PIN O1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.536 0.000 101.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.536 0.000 101.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.536 0.000 101.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.536 0.000 101.688 0.152 ;
    END
  END O1[54]

  PIN O1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.232 0.000 101.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.232 0.000 101.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.232 0.000 101.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.232 0.000 101.384 0.152 ;
    END
  END O1[53]

  PIN O1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.928 0.000 101.080 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.928 0.000 101.080 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.928 0.000 101.080 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.928 0.000 101.080 0.152 ;
    END
  END O1[52]

  PIN O1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.192 0.000 98.344 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.192 0.000 98.344 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.192 0.000 98.344 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.192 0.000 98.344 0.152 ;
    END
  END O1[59]

  PIN O1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.888 0.000 98.040 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.888 0.000 98.040 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.888 0.000 98.040 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.888 0.000 98.040 0.152 ;
    END
  END O1[58]

  PIN O1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.584 0.000 97.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.584 0.000 97.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.584 0.000 97.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.584 0.000 97.736 0.152 ;
    END
  END O1[57]

  PIN O1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.280 0.000 97.432 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.280 0.000 97.432 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.280 0.000 97.432 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.280 0.000 97.432 0.152 ;
    END
  END O1[56]

  PIN O1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.544 0.000 94.696 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.544 0.000 94.696 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.544 0.000 94.696 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.544 0.000 94.696 0.152 ;
    END
  END O1[63]

  PIN O1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 94.240 0.000 94.392 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 94.240 0.000 94.392 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 94.240 0.000 94.392 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 94.240 0.000 94.392 0.152 ;
    END
  END O1[62]

  PIN O1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.936 0.000 94.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.936 0.000 94.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.936 0.000 94.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.936 0.000 94.088 0.152 ;
    END
  END O1[61]

  PIN O1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.632 0.000 93.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.632 0.000 93.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.632 0.000 93.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.632 0.000 93.784 0.152 ;
    END
  END O1[60]

  PIN O1[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.896 0.000 91.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.896 0.000 91.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.896 0.000 91.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.896 0.000 91.048 0.152 ;
    END
  END O1[67]

  PIN O1[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.592 0.000 90.744 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.592 0.000 90.744 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.592 0.000 90.744 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.592 0.000 90.744 0.152 ;
    END
  END O1[66]

  PIN O1[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.288 0.000 90.440 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.288 0.000 90.440 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.288 0.000 90.440 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.288 0.000 90.440 0.152 ;
    END
  END O1[65]

  PIN O1[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.984 0.000 90.136 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.984 0.000 90.136 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.984 0.000 90.136 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.984 0.000 90.136 0.152 ;
    END
  END O1[64]

  PIN O1[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.248 0.000 87.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.248 0.000 87.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.248 0.000 87.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.248 0.000 87.400 0.152 ;
    END
  END O1[71]

  PIN O1[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.944 0.000 87.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.944 0.000 87.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.944 0.000 87.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.944 0.000 87.096 0.152 ;
    END
  END O1[70]

  PIN O1[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.640 0.000 86.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.640 0.000 86.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.640 0.000 86.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.640 0.000 86.792 0.152 ;
    END
  END O1[69]

  PIN O1[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.336 0.000 86.488 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.336 0.000 86.488 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.336 0.000 86.488 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.336 0.000 86.488 0.152 ;
    END
  END O1[68]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.576 64.904 161.728 65.056 ;
    END
    PORT
      LAYER M3 ;
        RECT 161.576 64.904 161.728 65.056 ;
    END
    PORT
      LAYER M4 ;
        RECT 161.576 64.904 161.728 65.056 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.576 64.904 161.728 65.056 ;
    END
  END A1[0]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.576 61.256 161.728 61.408 ;
    END
    PORT
      LAYER M3 ;
        RECT 161.576 61.256 161.728 61.408 ;
    END
    PORT
      LAYER M4 ;
        RECT 161.576 61.256 161.728 61.408 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.576 61.256 161.728 61.408 ;
    END
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.576 57.608 161.728 57.760 ;
    END
    PORT
      LAYER M3 ;
        RECT 161.576 57.608 161.728 57.760 ;
    END
    PORT
      LAYER M4 ;
        RECT 161.576 57.608 161.728 57.760 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.576 57.608 161.728 57.760 ;
    END
  END A1[2]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.576 53.960 161.728 54.112 ;
    END
    PORT
      LAYER M3 ;
        RECT 161.576 53.960 161.728 54.112 ;
    END
    PORT
      LAYER M4 ;
        RECT 161.576 53.960 161.728 54.112 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.576 53.960 161.728 54.112 ;
    END
  END A1[3]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.576 50.312 161.728 50.464 ;
    END
    PORT
      LAYER M3 ;
        RECT 161.576 50.312 161.728 50.464 ;
    END
    PORT
      LAYER M4 ;
        RECT 161.576 50.312 161.728 50.464 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.576 50.312 161.728 50.464 ;
    END
  END A1[4]

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.576 46.664 161.728 46.816 ;
    END
    PORT
      LAYER M3 ;
        RECT 161.576 46.664 161.728 46.816 ;
    END
    PORT
      LAYER M4 ;
        RECT 161.576 46.664 161.728 46.816 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.576 46.664 161.728 46.816 ;
    END
  END A1[5]

  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.576 43.016 161.728 43.168 ;
    END
    PORT
      LAYER M3 ;
        RECT 161.576 43.016 161.728 43.168 ;
    END
    PORT
      LAYER M4 ;
        RECT 161.576 43.016 161.728 43.168 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.576 43.016 161.728 43.168 ;
    END
  END A1[6]

  PIN A1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 161.576 39.368 161.728 39.520 ;
    END
    PORT
      LAYER M3 ;
        RECT 161.576 39.368 161.728 39.520 ;
    END
    PORT
      LAYER M4 ;
        RECT 161.576 39.368 161.728 39.520 ;
    END
    PORT
      LAYER M5 ;
        RECT 161.576 39.368 161.728 39.520 ;
    END
  END A1[7]

  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4.256 0.000 4.408 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 4.256 0.000 4.408 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 4.256 0.000 4.408 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 4.256 0.000 4.408 0.152 ;
    END
  END CE2

  PIN CSB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 6.992 0.000 7.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 6.992 0.000 7.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 6.992 0.000 7.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 6.992 0.000 7.144 0.152 ;
    END
  END CSB2

  PIN I2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.728 0.000 9.880 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 9.728 0.000 9.880 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 9.728 0.000 9.880 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 9.728 0.000 9.880 0.152 ;
    END
  END I2[0]

  PIN I2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.032 0.000 10.184 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.032 0.000 10.184 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.032 0.000 10.184 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.032 0.000 10.184 0.152 ;
    END
  END I2[1]

  PIN I2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.336 0.000 10.488 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.336 0.000 10.488 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.336 0.000 10.488 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.336 0.000 10.488 0.152 ;
    END
  END I2[2]

  PIN I2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 10.640 0.000 10.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 10.640 0.000 10.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 10.640 0.000 10.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 10.640 0.000 10.792 0.152 ;
    END
  END I2[3]

  PIN I2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.376 0.000 13.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.376 0.000 13.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.376 0.000 13.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.376 0.000 13.528 0.152 ;
    END
  END I2[4]

  PIN I2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.680 0.000 13.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.680 0.000 13.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.680 0.000 13.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.680 0.000 13.832 0.152 ;
    END
  END I2[5]

  PIN I2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.984 0.000 14.136 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 13.984 0.000 14.136 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 13.984 0.000 14.136 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 13.984 0.000 14.136 0.152 ;
    END
  END I2[6]

  PIN I2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.288 0.000 14.440 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 14.288 0.000 14.440 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 14.288 0.000 14.440 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 14.288 0.000 14.440 0.152 ;
    END
  END I2[7]

  PIN I2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.024 0.000 17.176 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.024 0.000 17.176 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.024 0.000 17.176 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.024 0.000 17.176 0.152 ;
    END
  END I2[8]

  PIN I2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.328 0.000 17.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.328 0.000 17.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.328 0.000 17.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.328 0.000 17.480 0.152 ;
    END
  END I2[9]

  PIN I2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.632 0.000 17.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.632 0.000 17.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.632 0.000 17.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.632 0.000 17.784 0.152 ;
    END
  END I2[10]

  PIN I2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 17.936 0.000 18.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 17.936 0.000 18.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 17.936 0.000 18.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 17.936 0.000 18.088 0.152 ;
    END
  END I2[11]

  PIN I2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.672 0.000 20.824 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.672 0.000 20.824 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.672 0.000 20.824 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.672 0.000 20.824 0.152 ;
    END
  END I2[12]

  PIN I2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.976 0.000 21.128 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.976 0.000 21.128 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.976 0.000 21.128 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.976 0.000 21.128 0.152 ;
    END
  END I2[13]

  PIN I2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.280 0.000 21.432 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.280 0.000 21.432 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.280 0.000 21.432 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.280 0.000 21.432 0.152 ;
    END
  END I2[14]

  PIN I2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.584 0.000 21.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.584 0.000 21.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.584 0.000 21.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.584 0.000 21.736 0.152 ;
    END
  END I2[15]

  PIN I2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.320 0.000 24.472 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.320 0.000 24.472 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.320 0.000 24.472 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.320 0.000 24.472 0.152 ;
    END
  END I2[16]

  PIN I2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.624 0.000 24.776 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.624 0.000 24.776 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.624 0.000 24.776 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.624 0.000 24.776 0.152 ;
    END
  END I2[17]

  PIN I2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.928 0.000 25.080 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.928 0.000 25.080 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.928 0.000 25.080 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.928 0.000 25.080 0.152 ;
    END
  END I2[18]

  PIN I2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.232 0.000 25.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.232 0.000 25.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.232 0.000 25.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.232 0.000 25.384 0.152 ;
    END
  END I2[19]

  PIN I2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
  END I2[20]

  PIN I2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.272 0.000 28.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.272 0.000 28.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.272 0.000 28.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.272 0.000 28.424 0.152 ;
    END
  END I2[21]

  PIN I2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.576 0.000 28.728 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.576 0.000 28.728 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.576 0.000 28.728 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.576 0.000 28.728 0.152 ;
    END
  END I2[22]

  PIN I2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.880 0.000 29.032 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 28.880 0.000 29.032 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 28.880 0.000 29.032 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 28.880 0.000 29.032 0.152 ;
    END
  END I2[23]

  PIN I2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.616 0.000 31.768 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.616 0.000 31.768 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.616 0.000 31.768 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.616 0.000 31.768 0.152 ;
    END
  END I2[24]

  PIN I2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
  END I2[25]

  PIN I2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.224 0.000 32.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.224 0.000 32.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.224 0.000 32.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.224 0.000 32.376 0.152 ;
    END
  END I2[26]

  PIN I2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.528 0.000 32.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.528 0.000 32.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.528 0.000 32.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.528 0.000 32.680 0.152 ;
    END
  END I2[27]

  PIN I2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.264 0.000 35.416 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.264 0.000 35.416 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.264 0.000 35.416 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.264 0.000 35.416 0.152 ;
    END
  END I2[28]

  PIN I2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.568 0.000 35.720 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.568 0.000 35.720 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.568 0.000 35.720 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.568 0.000 35.720 0.152 ;
    END
  END I2[29]

  PIN I2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.872 0.000 36.024 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.872 0.000 36.024 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.872 0.000 36.024 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.872 0.000 36.024 0.152 ;
    END
  END I2[30]

  PIN I2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.176 0.000 36.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.176 0.000 36.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.176 0.000 36.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.176 0.000 36.328 0.152 ;
    END
  END I2[31]

  PIN I2[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.912 0.000 39.064 0.152 ;
    END
  END I2[32]

  PIN I2[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.216 0.000 39.368 0.152 ;
    END
  END I2[33]

  PIN I2[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.520 0.000 39.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.520 0.000 39.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.520 0.000 39.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.520 0.000 39.672 0.152 ;
    END
  END I2[34]

  PIN I2[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.824 0.000 39.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.824 0.000 39.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.824 0.000 39.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.824 0.000 39.976 0.152 ;
    END
  END I2[35]

  PIN I2[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.560 0.000 42.712 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.560 0.000 42.712 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.560 0.000 42.712 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.560 0.000 42.712 0.152 ;
    END
  END I2[36]

  PIN I2[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.864 0.000 43.016 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.864 0.000 43.016 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.864 0.000 43.016 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.864 0.000 43.016 0.152 ;
    END
  END I2[37]

  PIN I2[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.168 0.000 43.320 0.152 ;
    END
  END I2[38]

  PIN I2[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 43.472 0.000 43.624 0.152 ;
    END
  END I2[39]

  PIN I2[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
  END I2[40]

  PIN I2[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.512 0.000 46.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.512 0.000 46.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.512 0.000 46.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.512 0.000 46.664 0.152 ;
    END
  END I2[41]

  PIN I2[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
  END I2[42]

  PIN I2[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
  END I2[43]

  PIN I2[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.856 0.000 50.008 0.152 ;
    END
  END I2[44]

  PIN I2[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.160 0.000 50.312 0.152 ;
    END
  END I2[45]

  PIN I2[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
  END I2[46]

  PIN I2[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.768 0.000 50.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.768 0.000 50.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.768 0.000 50.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.768 0.000 50.920 0.152 ;
    END
  END I2[47]

  PIN I2[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.504 0.000 53.656 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.504 0.000 53.656 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.504 0.000 53.656 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.504 0.000 53.656 0.152 ;
    END
  END I2[48]

  PIN I2[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.808 0.000 53.960 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.808 0.000 53.960 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.808 0.000 53.960 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.808 0.000 53.960 0.152 ;
    END
  END I2[49]

  PIN I2[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.112 0.000 54.264 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.112 0.000 54.264 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.112 0.000 54.264 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.112 0.000 54.264 0.152 ;
    END
  END I2[50]

  PIN I2[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.416 0.000 54.568 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.416 0.000 54.568 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.416 0.000 54.568 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.416 0.000 54.568 0.152 ;
    END
  END I2[51]

  PIN I2[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.152 0.000 57.304 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.152 0.000 57.304 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.152 0.000 57.304 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.152 0.000 57.304 0.152 ;
    END
  END I2[52]

  PIN I2[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.456 0.000 57.608 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.456 0.000 57.608 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.456 0.000 57.608 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.456 0.000 57.608 0.152 ;
    END
  END I2[53]

  PIN I2[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.760 0.000 57.912 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.760 0.000 57.912 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.760 0.000 57.912 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.760 0.000 57.912 0.152 ;
    END
  END I2[54]

  PIN I2[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.064 0.000 58.216 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.064 0.000 58.216 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.064 0.000 58.216 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.064 0.000 58.216 0.152 ;
    END
  END I2[55]

  PIN I2[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 60.800 0.000 60.952 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 60.800 0.000 60.952 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 60.800 0.000 60.952 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 60.800 0.000 60.952 0.152 ;
    END
  END I2[56]

  PIN I2[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.104 0.000 61.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.104 0.000 61.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.104 0.000 61.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.104 0.000 61.256 0.152 ;
    END
  END I2[57]

  PIN I2[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.408 0.000 61.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.408 0.000 61.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.408 0.000 61.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.408 0.000 61.560 0.152 ;
    END
  END I2[58]

  PIN I2[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.712 0.000 61.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.712 0.000 61.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.712 0.000 61.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.712 0.000 61.864 0.152 ;
    END
  END I2[59]

  PIN I2[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.448 0.000 64.600 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.448 0.000 64.600 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.448 0.000 64.600 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.448 0.000 64.600 0.152 ;
    END
  END I2[60]

  PIN I2[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.752 0.000 64.904 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.752 0.000 64.904 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.752 0.000 64.904 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.752 0.000 64.904 0.152 ;
    END
  END I2[61]

  PIN I2[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.056 0.000 65.208 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.056 0.000 65.208 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.056 0.000 65.208 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.056 0.000 65.208 0.152 ;
    END
  END I2[62]

  PIN I2[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.360 0.000 65.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.360 0.000 65.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.360 0.000 65.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.360 0.000 65.512 0.152 ;
    END
  END I2[63]

  PIN I2[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.096 0.000 68.248 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.096 0.000 68.248 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.096 0.000 68.248 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.096 0.000 68.248 0.152 ;
    END
  END I2[64]

  PIN I2[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.400 0.000 68.552 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.400 0.000 68.552 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.400 0.000 68.552 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.400 0.000 68.552 0.152 ;
    END
  END I2[65]

  PIN I2[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.704 0.000 68.856 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.704 0.000 68.856 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.704 0.000 68.856 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.704 0.000 68.856 0.152 ;
    END
  END I2[66]

  PIN I2[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.008 0.000 69.160 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.008 0.000 69.160 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.008 0.000 69.160 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.008 0.000 69.160 0.152 ;
    END
  END I2[67]

  PIN I2[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
  END I2[68]

  PIN I2[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.048 0.000 72.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.048 0.000 72.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.048 0.000 72.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.048 0.000 72.200 0.152 ;
    END
  END I2[69]

  PIN I2[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.352 0.000 72.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.352 0.000 72.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.352 0.000 72.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.352 0.000 72.504 0.152 ;
    END
  END I2[70]

  PIN I2[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.656 0.000 72.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.656 0.000 72.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.656 0.000 72.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.656 0.000 72.808 0.152 ;
    END
  END I2[71]

  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 64.904 0.152 65.056 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 64.904 0.152 65.056 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 64.904 0.152 65.056 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 64.904 0.152 65.056 ;
    END
  END A2[0]

  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 61.256 0.152 61.408 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 61.256 0.152 61.408 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 61.256 0.152 61.408 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 61.256 0.152 61.408 ;
    END
  END A2[1]

  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 57.608 0.152 57.760 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 57.608 0.152 57.760 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 57.608 0.152 57.760 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 57.608 0.152 57.760 ;
    END
  END A2[2]

  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 53.960 0.152 54.112 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 53.960 0.152 54.112 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 53.960 0.152 54.112 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 53.960 0.152 54.112 ;
    END
  END A2[3]

  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 50.312 0.152 50.464 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 50.312 0.152 50.464 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 50.312 0.152 50.464 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 50.312 0.152 50.464 ;
    END
  END A2[4]

  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 46.664 0.152 46.816 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 46.664 0.152 46.816 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 46.664 0.152 46.816 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 46.664 0.152 46.816 ;
    END
  END A2[5]

  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 43.016 0.152 43.168 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 43.016 0.152 43.168 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 43.016 0.152 43.168 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 43.016 0.152 43.168 ;
    END
  END A2[6]

  PIN A2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 39.368 0.152 39.520 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 39.368 0.152 39.520 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 39.368 0.152 39.520 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 39.368 0.152 39.520 ;
    END
  END A2[7]

  PIN WEB2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.000 18.544 0.152 18.696 ;
    END
    PORT
      LAYER M3 ;
        RECT 0.000 18.544 0.152 18.696 ;
    END
    PORT
      LAYER M4 ;
        RECT 0.000 18.544 0.152 18.696 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.000 18.544 0.152 18.696 ;
    END
  END WEB2

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 5.195 72.176 7.195 74.176 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.195 72.176 7.195 74.176 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.195 72.176 7.195 74.176 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M2 ;
        RECT 7.915 72.176 9.915 74.176 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.915 72.176 9.915 74.176 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.915 72.176 9.915 74.176 ;
    END
  END VSS

  OBS
    LAYER M2 ;
      RECT 157.776 0.000 161.728 0.304 ;
      RECT 155.040 0.000 157.320 0.304 ;
      RECT 152.304 0.000 154.584 0.304 ;
      RECT 149.568 0.000 151.848 0.304 ;
      RECT 145.920 0.000 148.200 0.304 ;
      RECT 142.272 0.000 144.552 0.304 ;
      RECT 138.624 0.000 140.904 0.304 ;
      RECT 134.976 0.000 137.256 0.304 ;
      RECT 131.328 0.000 133.608 0.304 ;
      RECT 127.680 0.000 129.960 0.304 ;
      RECT 124.032 0.000 126.312 0.304 ;
      RECT 120.384 0.000 122.664 0.304 ;
      RECT 116.736 0.000 119.016 0.304 ;
      RECT 113.088 0.000 115.368 0.304 ;
      RECT 109.440 0.000 111.720 0.304 ;
      RECT 105.792 0.000 108.072 0.304 ;
      RECT 102.144 0.000 104.424 0.304 ;
      RECT 98.496 0.000 100.776 0.304 ;
      RECT 94.848 0.000 97.128 0.304 ;
      RECT 91.200 0.000 93.480 0.304 ;
      RECT 87.552 0.000 89.832 0.304 ;
      RECT 161.424 65.208 161.728 72.024 ;
      RECT 161.424 61.560 161.728 64.752 ;
      RECT 161.424 57.912 161.728 61.104 ;
      RECT 161.424 54.264 161.728 57.456 ;
      RECT 161.424 50.616 161.728 53.808 ;
      RECT 161.424 46.968 161.728 50.160 ;
      RECT 161.424 43.320 161.728 46.512 ;
      RECT 161.424 39.672 161.728 42.864 ;
      RECT 161.424 18.848 161.728 39.216 ;
      RECT 161.424 0.304 161.728 18.392 ;
      RECT 0.000 0.000 4.104 0.304 ;
      RECT 4.560 0.000 6.840 0.304 ;
      RECT 7.296 0.000 9.576 0.304 ;
      RECT 10.944 0.000 13.224 0.304 ;
      RECT 14.592 0.000 16.872 0.304 ;
      RECT 18.240 0.000 20.520 0.304 ;
      RECT 21.888 0.000 24.168 0.304 ;
      RECT 25.536 0.000 27.816 0.304 ;
      RECT 29.184 0.000 31.464 0.304 ;
      RECT 32.832 0.000 35.112 0.304 ;
      RECT 36.480 0.000 38.760 0.304 ;
      RECT 40.128 0.000 42.408 0.304 ;
      RECT 43.776 0.000 46.056 0.304 ;
      RECT 47.424 0.000 49.704 0.304 ;
      RECT 51.072 0.000 53.352 0.304 ;
      RECT 54.720 0.000 57.000 0.304 ;
      RECT 58.368 0.000 60.648 0.304 ;
      RECT 62.016 0.000 64.296 0.304 ;
      RECT 65.664 0.000 67.944 0.304 ;
      RECT 69.312 0.000 71.592 0.304 ;
      RECT 72.960 0.000 86.184 0.304 ;
      RECT 0.000 65.208 0.304 72.024 ;
      RECT 0.000 61.560 0.304 64.752 ;
      RECT 0.000 57.912 0.304 61.104 ;
      RECT 0.000 54.264 0.304 57.456 ;
      RECT 0.000 50.616 0.304 53.808 ;
      RECT 0.000 46.968 0.304 50.160 ;
      RECT 0.000 43.320 0.304 46.512 ;
      RECT 0.000 39.672 0.304 42.864 ;
      RECT 0.000 18.848 0.304 39.216 ;
      RECT 0.000 0.304 0.304 18.392 ;
      RECT 0.000 72.024 5.043 74.176 ;
      RECT 7.355 72.024 7.763 74.176 ;
      RECT 10.067 72.024 161.728 74.176 ;
      RECT 0.304 0.304 161.424 72.024 ;
    LAYER M3 ;
      RECT 157.776 0.000 161.728 0.304 ;
      RECT 155.040 0.000 157.320 0.304 ;
      RECT 152.304 0.000 154.584 0.304 ;
      RECT 149.568 0.000 151.848 0.304 ;
      RECT 145.920 0.000 148.200 0.304 ;
      RECT 142.272 0.000 144.552 0.304 ;
      RECT 138.624 0.000 140.904 0.304 ;
      RECT 134.976 0.000 137.256 0.304 ;
      RECT 131.328 0.000 133.608 0.304 ;
      RECT 127.680 0.000 129.960 0.304 ;
      RECT 124.032 0.000 126.312 0.304 ;
      RECT 120.384 0.000 122.664 0.304 ;
      RECT 116.736 0.000 119.016 0.304 ;
      RECT 113.088 0.000 115.368 0.304 ;
      RECT 109.440 0.000 111.720 0.304 ;
      RECT 105.792 0.000 108.072 0.304 ;
      RECT 102.144 0.000 104.424 0.304 ;
      RECT 98.496 0.000 100.776 0.304 ;
      RECT 94.848 0.000 97.128 0.304 ;
      RECT 91.200 0.000 93.480 0.304 ;
      RECT 87.552 0.000 89.832 0.304 ;
      RECT 161.424 65.208 161.728 72.024 ;
      RECT 161.424 61.560 161.728 64.752 ;
      RECT 161.424 57.912 161.728 61.104 ;
      RECT 161.424 54.264 161.728 57.456 ;
      RECT 161.424 50.616 161.728 53.808 ;
      RECT 161.424 46.968 161.728 50.160 ;
      RECT 161.424 43.320 161.728 46.512 ;
      RECT 161.424 39.672 161.728 42.864 ;
      RECT 161.424 18.848 161.728 39.216 ;
      RECT 161.424 0.304 161.728 18.392 ;
      RECT 0.000 0.000 4.104 0.304 ;
      RECT 4.560 0.000 6.840 0.304 ;
      RECT 7.296 0.000 9.576 0.304 ;
      RECT 10.944 0.000 13.224 0.304 ;
      RECT 14.592 0.000 16.872 0.304 ;
      RECT 18.240 0.000 20.520 0.304 ;
      RECT 21.888 0.000 24.168 0.304 ;
      RECT 25.536 0.000 27.816 0.304 ;
      RECT 29.184 0.000 31.464 0.304 ;
      RECT 32.832 0.000 35.112 0.304 ;
      RECT 36.480 0.000 38.760 0.304 ;
      RECT 40.128 0.000 42.408 0.304 ;
      RECT 43.776 0.000 46.056 0.304 ;
      RECT 47.424 0.000 49.704 0.304 ;
      RECT 51.072 0.000 53.352 0.304 ;
      RECT 54.720 0.000 57.000 0.304 ;
      RECT 58.368 0.000 60.648 0.304 ;
      RECT 62.016 0.000 64.296 0.304 ;
      RECT 65.664 0.000 67.944 0.304 ;
      RECT 69.312 0.000 71.592 0.304 ;
      RECT 72.960 0.000 86.184 0.304 ;
      RECT 0.000 65.208 0.304 72.024 ;
      RECT 0.000 61.560 0.304 64.752 ;
      RECT 0.000 57.912 0.304 61.104 ;
      RECT 0.000 54.264 0.304 57.456 ;
      RECT 0.000 50.616 0.304 53.808 ;
      RECT 0.000 46.968 0.304 50.160 ;
      RECT 0.000 43.320 0.304 46.512 ;
      RECT 0.000 39.672 0.304 42.864 ;
      RECT 0.000 18.848 0.304 39.216 ;
      RECT 0.000 0.304 0.304 18.392 ;
      RECT 0.000 72.024 5.043 74.176 ;
      RECT 7.355 72.024 7.763 74.176 ;
      RECT 10.067 72.024 161.728 74.176 ;
      RECT 0.304 0.304 161.424 72.024 ;
    LAYER M4 ;
      RECT 157.776 0.000 161.728 0.304 ;
      RECT 155.040 0.000 157.320 0.304 ;
      RECT 152.304 0.000 154.584 0.304 ;
      RECT 149.568 0.000 151.848 0.304 ;
      RECT 145.920 0.000 148.200 0.304 ;
      RECT 142.272 0.000 144.552 0.304 ;
      RECT 138.624 0.000 140.904 0.304 ;
      RECT 134.976 0.000 137.256 0.304 ;
      RECT 131.328 0.000 133.608 0.304 ;
      RECT 127.680 0.000 129.960 0.304 ;
      RECT 124.032 0.000 126.312 0.304 ;
      RECT 120.384 0.000 122.664 0.304 ;
      RECT 116.736 0.000 119.016 0.304 ;
      RECT 113.088 0.000 115.368 0.304 ;
      RECT 109.440 0.000 111.720 0.304 ;
      RECT 105.792 0.000 108.072 0.304 ;
      RECT 102.144 0.000 104.424 0.304 ;
      RECT 98.496 0.000 100.776 0.304 ;
      RECT 94.848 0.000 97.128 0.304 ;
      RECT 91.200 0.000 93.480 0.304 ;
      RECT 87.552 0.000 89.832 0.304 ;
      RECT 161.424 65.208 161.728 72.024 ;
      RECT 161.424 61.560 161.728 64.752 ;
      RECT 161.424 57.912 161.728 61.104 ;
      RECT 161.424 54.264 161.728 57.456 ;
      RECT 161.424 50.616 161.728 53.808 ;
      RECT 161.424 46.968 161.728 50.160 ;
      RECT 161.424 43.320 161.728 46.512 ;
      RECT 161.424 39.672 161.728 42.864 ;
      RECT 161.424 18.848 161.728 39.216 ;
      RECT 161.424 0.304 161.728 18.392 ;
      RECT 0.000 0.000 4.104 0.304 ;
      RECT 4.560 0.000 6.840 0.304 ;
      RECT 7.296 0.000 9.576 0.304 ;
      RECT 10.944 0.000 13.224 0.304 ;
      RECT 14.592 0.000 16.872 0.304 ;
      RECT 18.240 0.000 20.520 0.304 ;
      RECT 21.888 0.000 24.168 0.304 ;
      RECT 25.536 0.000 27.816 0.304 ;
      RECT 29.184 0.000 31.464 0.304 ;
      RECT 32.832 0.000 35.112 0.304 ;
      RECT 36.480 0.000 38.760 0.304 ;
      RECT 40.128 0.000 42.408 0.304 ;
      RECT 43.776 0.000 46.056 0.304 ;
      RECT 47.424 0.000 49.704 0.304 ;
      RECT 51.072 0.000 53.352 0.304 ;
      RECT 54.720 0.000 57.000 0.304 ;
      RECT 58.368 0.000 60.648 0.304 ;
      RECT 62.016 0.000 64.296 0.304 ;
      RECT 65.664 0.000 67.944 0.304 ;
      RECT 69.312 0.000 71.592 0.304 ;
      RECT 72.960 0.000 86.184 0.304 ;
      RECT 0.000 65.208 0.304 72.024 ;
      RECT 0.000 61.560 0.304 64.752 ;
      RECT 0.000 57.912 0.304 61.104 ;
      RECT 0.000 54.264 0.304 57.456 ;
      RECT 0.000 50.616 0.304 53.808 ;
      RECT 0.000 46.968 0.304 50.160 ;
      RECT 0.000 43.320 0.304 46.512 ;
      RECT 0.000 39.672 0.304 42.864 ;
      RECT 0.000 18.848 0.304 39.216 ;
      RECT 0.000 0.304 0.304 18.392 ;
      RECT 0.000 72.024 5.043 74.176 ;
      RECT 7.355 72.024 7.763 74.176 ;
      RECT 10.067 72.024 161.728 74.176 ;
      RECT 0.304 0.304 161.424 72.024 ;
    LAYER M5 ;
      RECT 157.776 0.000 161.728 0.304 ;
      RECT 155.040 0.000 157.320 0.304 ;
      RECT 152.304 0.000 154.584 0.304 ;
      RECT 149.568 0.000 151.848 0.304 ;
      RECT 145.920 0.000 148.200 0.304 ;
      RECT 142.272 0.000 144.552 0.304 ;
      RECT 138.624 0.000 140.904 0.304 ;
      RECT 134.976 0.000 137.256 0.304 ;
      RECT 131.328 0.000 133.608 0.304 ;
      RECT 127.680 0.000 129.960 0.304 ;
      RECT 124.032 0.000 126.312 0.304 ;
      RECT 120.384 0.000 122.664 0.304 ;
      RECT 116.736 0.000 119.016 0.304 ;
      RECT 113.088 0.000 115.368 0.304 ;
      RECT 109.440 0.000 111.720 0.304 ;
      RECT 105.792 0.000 108.072 0.304 ;
      RECT 102.144 0.000 104.424 0.304 ;
      RECT 98.496 0.000 100.776 0.304 ;
      RECT 94.848 0.000 97.128 0.304 ;
      RECT 91.200 0.000 93.480 0.304 ;
      RECT 87.552 0.000 89.832 0.304 ;
      RECT 161.424 65.208 161.728 72.024 ;
      RECT 161.424 61.560 161.728 64.752 ;
      RECT 161.424 57.912 161.728 61.104 ;
      RECT 161.424 54.264 161.728 57.456 ;
      RECT 161.424 50.616 161.728 53.808 ;
      RECT 161.424 46.968 161.728 50.160 ;
      RECT 161.424 43.320 161.728 46.512 ;
      RECT 161.424 39.672 161.728 42.864 ;
      RECT 161.424 18.848 161.728 39.216 ;
      RECT 161.424 0.304 161.728 18.392 ;
      RECT 0.000 0.000 4.104 0.304 ;
      RECT 4.560 0.000 6.840 0.304 ;
      RECT 7.296 0.000 9.576 0.304 ;
      RECT 10.944 0.000 13.224 0.304 ;
      RECT 14.592 0.000 16.872 0.304 ;
      RECT 18.240 0.000 20.520 0.304 ;
      RECT 21.888 0.000 24.168 0.304 ;
      RECT 25.536 0.000 27.816 0.304 ;
      RECT 29.184 0.000 31.464 0.304 ;
      RECT 32.832 0.000 35.112 0.304 ;
      RECT 36.480 0.000 38.760 0.304 ;
      RECT 40.128 0.000 42.408 0.304 ;
      RECT 43.776 0.000 46.056 0.304 ;
      RECT 47.424 0.000 49.704 0.304 ;
      RECT 51.072 0.000 53.352 0.304 ;
      RECT 54.720 0.000 57.000 0.304 ;
      RECT 58.368 0.000 60.648 0.304 ;
      RECT 62.016 0.000 64.296 0.304 ;
      RECT 65.664 0.000 67.944 0.304 ;
      RECT 69.312 0.000 71.592 0.304 ;
      RECT 72.960 0.000 86.184 0.304 ;
      RECT 0.000 65.208 0.304 72.024 ;
      RECT 0.000 61.560 0.304 64.752 ;
      RECT 0.000 57.912 0.304 61.104 ;
      RECT 0.000 54.264 0.304 57.456 ;
      RECT 0.000 50.616 0.304 53.808 ;
      RECT 0.000 46.968 0.304 50.160 ;
      RECT 0.000 43.320 0.304 46.512 ;
      RECT 0.000 39.672 0.304 42.864 ;
      RECT 0.000 18.848 0.304 39.216 ;
      RECT 0.000 0.304 0.304 18.392 ;
      RECT 0.000 72.024 5.043 74.176 ;
      RECT 7.355 72.024 7.763 74.176 ;
      RECT 10.067 72.024 161.728 74.176 ;
      RECT 0.304 0.304 161.424 72.024 ;
  END

END sram8t256x72

END LIBRARY
