VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram6t512x128
  CLASS BLOCK ;
  SOURCE USER ;
  ORIGIN 0 0 ;
  SIZE 177.536 BY 97.280 ;
  SYMMETRY X Y R90 ;

  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.296 0.000 159.448 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 159.296 0.000 159.448 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 159.296 0.000 159.448 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 159.296 0.000 159.448 0.152 ;
    END
  END CE1

  PIN CSB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 158.080 0.000 158.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 158.080 0.000 158.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 158.080 0.000 158.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 158.080 0.000 158.232 0.152 ;
    END
  END CSB1

  PIN OEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 156.864 0.000 157.016 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 156.864 0.000 157.016 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 156.864 0.000 157.016 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 156.864 0.000 157.016 0.152 ;
    END
  END OEB1

  PIN O1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.648 0.000 155.800 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 155.648 0.000 155.800 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 155.648 0.000 155.800 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 155.648 0.000 155.800 0.152 ;
    END
  END O1[3]

  PIN O1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.344 0.000 155.496 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 155.344 0.000 155.496 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 155.344 0.000 155.496 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 155.344 0.000 155.496 0.152 ;
    END
  END O1[2]

  PIN O1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.040 0.000 155.192 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 155.040 0.000 155.192 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 155.040 0.000 155.192 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 155.040 0.000 155.192 0.152 ;
    END
  END O1[1]

  PIN O1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.736 0.000 154.888 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 154.736 0.000 154.888 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 154.736 0.000 154.888 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 154.736 0.000 154.888 0.152 ;
    END
  END O1[0]

  PIN I1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.520 0.000 153.672 0.152 ;
    END
  END I1[0]

  PIN I1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 153.216 0.000 153.368 0.152 ;
    END
  END I1[1]

  PIN I1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.912 0.000 153.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 152.912 0.000 153.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 152.912 0.000 153.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 152.912 0.000 153.064 0.152 ;
    END
  END I1[2]

  PIN I1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.608 0.000 152.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 152.608 0.000 152.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 152.608 0.000 152.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 152.608 0.000 152.760 0.152 ;
    END
  END I1[3]

  PIN O1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 151.392 0.000 151.544 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 151.392 0.000 151.544 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 151.392 0.000 151.544 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 151.392 0.000 151.544 0.152 ;
    END
  END O1[7]

  PIN O1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 151.088 0.000 151.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 151.088 0.000 151.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 151.088 0.000 151.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 151.088 0.000 151.240 0.152 ;
    END
  END O1[6]

  PIN O1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.784 0.000 150.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.784 0.000 150.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.784 0.000 150.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 150.784 0.000 150.936 0.152 ;
    END
  END O1[5]

  PIN O1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 150.480 0.000 150.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 150.480 0.000 150.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.480 0.000 150.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 150.480 0.000 150.632 0.152 ;
    END
  END O1[4]

  PIN I1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.264 0.000 149.416 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 149.264 0.000 149.416 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 149.264 0.000 149.416 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 149.264 0.000 149.416 0.152 ;
    END
  END I1[4]

  PIN I1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.960 0.000 149.112 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.960 0.000 149.112 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.960 0.000 149.112 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.960 0.000 149.112 0.152 ;
    END
  END I1[5]

  PIN I1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.656 0.000 148.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.656 0.000 148.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.656 0.000 148.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.656 0.000 148.808 0.152 ;
    END
  END I1[6]

  PIN I1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.352 0.000 148.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 148.352 0.000 148.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 148.352 0.000 148.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 148.352 0.000 148.504 0.152 ;
    END
  END I1[7]

  PIN O1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.136 0.000 147.288 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 147.136 0.000 147.288 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 147.136 0.000 147.288 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 147.136 0.000 147.288 0.152 ;
    END
  END O1[11]

  PIN O1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.832 0.000 146.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 146.832 0.000 146.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 146.832 0.000 146.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.832 0.000 146.984 0.152 ;
    END
  END O1[10]

  PIN O1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.528 0.000 146.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 146.528 0.000 146.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 146.528 0.000 146.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.528 0.000 146.680 0.152 ;
    END
  END O1[9]

  PIN O1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.224 0.000 146.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 146.224 0.000 146.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 146.224 0.000 146.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 146.224 0.000 146.376 0.152 ;
    END
  END O1[8]

  PIN I1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.008 0.000 145.160 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 145.008 0.000 145.160 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 145.008 0.000 145.160 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 145.008 0.000 145.160 0.152 ;
    END
  END I1[8]

  PIN I1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.704 0.000 144.856 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 144.704 0.000 144.856 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 144.704 0.000 144.856 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 144.704 0.000 144.856 0.152 ;
    END
  END I1[9]

  PIN I1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.400 0.000 144.552 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 144.400 0.000 144.552 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 144.400 0.000 144.552 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 144.400 0.000 144.552 0.152 ;
    END
  END I1[10]

  PIN I1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.096 0.000 144.248 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 144.096 0.000 144.248 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 144.096 0.000 144.248 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 144.096 0.000 144.248 0.152 ;
    END
  END I1[11]

  PIN O1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.880 0.000 143.032 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 142.880 0.000 143.032 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 142.880 0.000 143.032 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 142.880 0.000 143.032 0.152 ;
    END
  END O1[15]

  PIN O1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.576 0.000 142.728 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 142.576 0.000 142.728 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 142.576 0.000 142.728 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 142.576 0.000 142.728 0.152 ;
    END
  END O1[14]

  PIN O1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 142.272 0.000 142.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 142.272 0.000 142.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 142.272 0.000 142.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 142.272 0.000 142.424 0.152 ;
    END
  END O1[13]

  PIN O1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.968 0.000 142.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 141.968 0.000 142.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 141.968 0.000 142.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 141.968 0.000 142.120 0.152 ;
    END
  END O1[12]

  PIN I1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.752 0.000 140.904 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 140.752 0.000 140.904 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 140.752 0.000 140.904 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 140.752 0.000 140.904 0.152 ;
    END
  END I1[12]

  PIN I1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.448 0.000 140.600 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 140.448 0.000 140.600 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 140.448 0.000 140.600 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 140.448 0.000 140.600 0.152 ;
    END
  END I1[13]

  PIN I1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.144 0.000 140.296 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 140.144 0.000 140.296 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 140.144 0.000 140.296 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 140.144 0.000 140.296 0.152 ;
    END
  END I1[14]

  PIN I1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.840 0.000 139.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 139.840 0.000 139.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 139.840 0.000 139.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 139.840 0.000 139.992 0.152 ;
    END
  END I1[15]

  PIN O1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.624 0.000 138.776 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 138.624 0.000 138.776 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 138.624 0.000 138.776 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 138.624 0.000 138.776 0.152 ;
    END
  END O1[19]

  PIN O1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.320 0.000 138.472 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 138.320 0.000 138.472 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 138.320 0.000 138.472 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 138.320 0.000 138.472 0.152 ;
    END
  END O1[18]

  PIN O1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.016 0.000 138.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 138.016 0.000 138.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 138.016 0.000 138.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 138.016 0.000 138.168 0.152 ;
    END
  END O1[17]

  PIN O1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 137.712 0.000 137.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 137.712 0.000 137.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 137.712 0.000 137.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 137.712 0.000 137.864 0.152 ;
    END
  END O1[16]

  PIN I1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.496 0.000 136.648 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 136.496 0.000 136.648 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 136.496 0.000 136.648 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 136.496 0.000 136.648 0.152 ;
    END
  END I1[16]

  PIN I1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.192 0.000 136.344 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 136.192 0.000 136.344 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 136.192 0.000 136.344 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 136.192 0.000 136.344 0.152 ;
    END
  END I1[17]

  PIN I1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.888 0.000 136.040 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 135.888 0.000 136.040 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 135.888 0.000 136.040 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 135.888 0.000 136.040 0.152 ;
    END
  END I1[18]

  PIN I1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.584 0.000 135.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 135.584 0.000 135.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 135.584 0.000 135.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 135.584 0.000 135.736 0.152 ;
    END
  END I1[19]

  PIN O1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.368 0.000 134.520 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 134.368 0.000 134.520 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 134.368 0.000 134.520 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.368 0.000 134.520 0.152 ;
    END
  END O1[23]

  PIN O1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.064 0.000 134.216 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 134.064 0.000 134.216 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 134.064 0.000 134.216 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 134.064 0.000 134.216 0.152 ;
    END
  END O1[22]

  PIN O1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.760 0.000 133.912 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 133.760 0.000 133.912 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 133.760 0.000 133.912 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 133.760 0.000 133.912 0.152 ;
    END
  END O1[21]

  PIN O1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.456 0.000 133.608 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 133.456 0.000 133.608 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 133.456 0.000 133.608 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 133.456 0.000 133.608 0.152 ;
    END
  END O1[20]

  PIN I1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.240 0.000 132.392 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 132.240 0.000 132.392 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 132.240 0.000 132.392 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 132.240 0.000 132.392 0.152 ;
    END
  END I1[20]

  PIN I1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.936 0.000 132.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.936 0.000 132.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.936 0.000 132.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.936 0.000 132.088 0.152 ;
    END
  END I1[21]

  PIN I1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.632 0.000 131.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.632 0.000 131.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.632 0.000 131.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.632 0.000 131.784 0.152 ;
    END
  END I1[22]

  PIN I1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.328 0.000 131.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 131.328 0.000 131.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 131.328 0.000 131.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 131.328 0.000 131.480 0.152 ;
    END
  END I1[23]

  PIN O1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.112 0.000 130.264 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 130.112 0.000 130.264 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 130.112 0.000 130.264 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 130.112 0.000 130.264 0.152 ;
    END
  END O1[27]

  PIN O1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.808 0.000 129.960 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 129.808 0.000 129.960 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 129.808 0.000 129.960 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.808 0.000 129.960 0.152 ;
    END
  END O1[26]

  PIN O1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.504 0.000 129.656 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 129.504 0.000 129.656 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 129.504 0.000 129.656 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.504 0.000 129.656 0.152 ;
    END
  END O1[25]

  PIN O1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 129.200 0.000 129.352 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 129.200 0.000 129.352 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 129.200 0.000 129.352 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 129.200 0.000 129.352 0.152 ;
    END
  END O1[24]

  PIN I1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.984 0.000 128.136 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 127.984 0.000 128.136 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 127.984 0.000 128.136 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.984 0.000 128.136 0.152 ;
    END
  END I1[24]

  PIN I1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.680 0.000 127.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 127.680 0.000 127.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 127.680 0.000 127.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.680 0.000 127.832 0.152 ;
    END
  END I1[25]

  PIN I1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.376 0.000 127.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 127.376 0.000 127.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 127.376 0.000 127.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.376 0.000 127.528 0.152 ;
    END
  END I1[26]

  PIN I1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.072 0.000 127.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 127.072 0.000 127.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 127.072 0.000 127.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 127.072 0.000 127.224 0.152 ;
    END
  END I1[27]

  PIN O1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.856 0.000 126.008 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 125.856 0.000 126.008 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 125.856 0.000 126.008 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.856 0.000 126.008 0.152 ;
    END
  END O1[31]

  PIN O1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.552 0.000 125.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 125.552 0.000 125.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 125.552 0.000 125.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.552 0.000 125.704 0.152 ;
    END
  END O1[30]

  PIN O1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.248 0.000 125.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 125.248 0.000 125.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 125.248 0.000 125.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 125.248 0.000 125.400 0.152 ;
    END
  END O1[29]

  PIN O1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.944 0.000 125.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 124.944 0.000 125.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 124.944 0.000 125.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 124.944 0.000 125.096 0.152 ;
    END
  END O1[28]

  PIN I1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.728 0.000 123.880 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 123.728 0.000 123.880 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 123.728 0.000 123.880 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.728 0.000 123.880 0.152 ;
    END
  END I1[28]

  PIN I1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.424 0.000 123.576 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 123.424 0.000 123.576 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 123.424 0.000 123.576 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.424 0.000 123.576 0.152 ;
    END
  END I1[29]

  PIN I1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.120 0.000 123.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 123.120 0.000 123.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 123.120 0.000 123.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 123.120 0.000 123.272 0.152 ;
    END
  END I1[30]

  PIN I1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.816 0.000 122.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 122.816 0.000 122.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 122.816 0.000 122.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 122.816 0.000 122.968 0.152 ;
    END
  END I1[31]

  PIN O1[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.600 0.000 121.752 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 121.600 0.000 121.752 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 121.600 0.000 121.752 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.600 0.000 121.752 0.152 ;
    END
  END O1[35]

  PIN O1[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 121.296 0.000 121.448 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 121.296 0.000 121.448 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 121.296 0.000 121.448 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 121.296 0.000 121.448 0.152 ;
    END
  END O1[34]

  PIN O1[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.992 0.000 121.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.992 0.000 121.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.992 0.000 121.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.992 0.000 121.144 0.152 ;
    END
  END O1[33]

  PIN O1[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.688 0.000 120.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 120.688 0.000 120.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 120.688 0.000 120.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 120.688 0.000 120.840 0.152 ;
    END
  END O1[32]

  PIN I1[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.472 0.000 119.624 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 119.472 0.000 119.624 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 119.472 0.000 119.624 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.472 0.000 119.624 0.152 ;
    END
  END I1[32]

  PIN I1[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.168 0.000 119.320 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 119.168 0.000 119.320 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 119.168 0.000 119.320 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 119.168 0.000 119.320 0.152 ;
    END
  END I1[33]

  PIN I1[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.864 0.000 119.016 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 118.864 0.000 119.016 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 118.864 0.000 119.016 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.864 0.000 119.016 0.152 ;
    END
  END I1[34]

  PIN I1[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 118.560 0.000 118.712 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 118.560 0.000 118.712 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 118.560 0.000 118.712 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 118.560 0.000 118.712 0.152 ;
    END
  END I1[35]

  PIN O1[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.344 0.000 117.496 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 117.344 0.000 117.496 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 117.344 0.000 117.496 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.344 0.000 117.496 0.152 ;
    END
  END O1[39]

  PIN O1[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.040 0.000 117.192 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 117.040 0.000 117.192 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 117.040 0.000 117.192 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 117.040 0.000 117.192 0.152 ;
    END
  END O1[38]

  PIN O1[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.736 0.000 116.888 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 116.736 0.000 116.888 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 116.736 0.000 116.888 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.736 0.000 116.888 0.152 ;
    END
  END O1[37]

  PIN O1[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 116.432 0.000 116.584 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 116.432 0.000 116.584 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 116.432 0.000 116.584 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 116.432 0.000 116.584 0.152 ;
    END
  END O1[36]

  PIN I1[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.216 0.000 115.368 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 115.216 0.000 115.368 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 115.216 0.000 115.368 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 115.216 0.000 115.368 0.152 ;
    END
  END I1[36]

  PIN I1[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.912 0.000 115.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 114.912 0.000 115.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 114.912 0.000 115.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.912 0.000 115.064 0.152 ;
    END
  END I1[37]

  PIN I1[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.608 0.000 114.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 114.608 0.000 114.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 114.608 0.000 114.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.608 0.000 114.760 0.152 ;
    END
  END I1[38]

  PIN I1[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.304 0.000 114.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 114.304 0.000 114.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 114.304 0.000 114.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 114.304 0.000 114.456 0.152 ;
    END
  END I1[39]

  PIN O1[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 113.088 0.000 113.240 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 113.088 0.000 113.240 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 113.088 0.000 113.240 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 113.088 0.000 113.240 0.152 ;
    END
  END O1[43]

  PIN O1[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.784 0.000 112.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 112.784 0.000 112.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.784 0.000 112.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.784 0.000 112.936 0.152 ;
    END
  END O1[42]

  PIN O1[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.480 0.000 112.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 112.480 0.000 112.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.480 0.000 112.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.480 0.000 112.632 0.152 ;
    END
  END O1[41]

  PIN O1[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.176 0.000 112.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 112.176 0.000 112.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 112.176 0.000 112.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 112.176 0.000 112.328 0.152 ;
    END
  END O1[40]

  PIN I1[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.960 0.000 111.112 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.960 0.000 111.112 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.960 0.000 111.112 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.960 0.000 111.112 0.152 ;
    END
  END I1[40]

  PIN I1[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.656 0.000 110.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.656 0.000 110.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.656 0.000 110.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.656 0.000 110.808 0.152 ;
    END
  END I1[41]

  PIN I1[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.352 0.000 110.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.352 0.000 110.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.352 0.000 110.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.352 0.000 110.504 0.152 ;
    END
  END I1[42]

  PIN I1[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 110.048 0.000 110.200 0.152 ;
    END
  END I1[43]

  PIN O1[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.832 0.000 108.984 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.832 0.000 108.984 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.832 0.000 108.984 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.832 0.000 108.984 0.152 ;
    END
  END O1[47]

  PIN O1[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.528 0.000 108.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.528 0.000 108.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.528 0.000 108.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.528 0.000 108.680 0.152 ;
    END
  END O1[46]

  PIN O1[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 108.224 0.000 108.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 108.224 0.000 108.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 108.224 0.000 108.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 108.224 0.000 108.376 0.152 ;
    END
  END O1[45]

  PIN O1[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.920 0.000 108.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 107.920 0.000 108.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 107.920 0.000 108.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 107.920 0.000 108.072 0.152 ;
    END
  END O1[44]

  PIN I1[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.704 0.000 106.856 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 106.704 0.000 106.856 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 106.704 0.000 106.856 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.704 0.000 106.856 0.152 ;
    END
  END I1[44]

  PIN I1[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.400 0.000 106.552 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 106.400 0.000 106.552 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 106.400 0.000 106.552 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.400 0.000 106.552 0.152 ;
    END
  END I1[45]

  PIN I1[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.096 0.000 106.248 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 106.096 0.000 106.248 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 106.096 0.000 106.248 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 106.096 0.000 106.248 0.152 ;
    END
  END I1[46]

  PIN I1[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.792 0.000 105.944 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 105.792 0.000 105.944 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 105.792 0.000 105.944 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 105.792 0.000 105.944 0.152 ;
    END
  END I1[47]

  PIN O1[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.576 0.000 104.728 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.576 0.000 104.728 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.576 0.000 104.728 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.576 0.000 104.728 0.152 ;
    END
  END O1[51]

  PIN O1[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.272 0.000 104.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 104.272 0.000 104.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 104.272 0.000 104.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 104.272 0.000 104.424 0.152 ;
    END
  END O1[50]

  PIN O1[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.968 0.000 104.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.968 0.000 104.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.968 0.000 104.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.968 0.000 104.120 0.152 ;
    END
  END O1[49]

  PIN O1[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.664 0.000 103.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 103.664 0.000 103.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 103.664 0.000 103.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 103.664 0.000 103.816 0.152 ;
    END
  END O1[48]

  PIN I1[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.448 0.000 102.600 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.448 0.000 102.600 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.448 0.000 102.600 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.448 0.000 102.600 0.152 ;
    END
  END I1[48]

  PIN I1[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 102.144 0.000 102.296 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 102.144 0.000 102.296 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 102.144 0.000 102.296 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 102.144 0.000 102.296 0.152 ;
    END
  END I1[49]

  PIN I1[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.840 0.000 101.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.840 0.000 101.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.840 0.000 101.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.840 0.000 101.992 0.152 ;
    END
  END I1[50]

  PIN I1[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.536 0.000 101.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 101.536 0.000 101.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 101.536 0.000 101.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 101.536 0.000 101.688 0.152 ;
    END
  END I1[51]

  PIN O1[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.320 0.000 100.472 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.320 0.000 100.472 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.320 0.000 100.472 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.320 0.000 100.472 0.152 ;
    END
  END O1[55]

  PIN O1[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.016 0.000 100.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 100.016 0.000 100.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 100.016 0.000 100.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 100.016 0.000 100.168 0.152 ;
    END
  END O1[54]

  PIN O1[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.712 0.000 99.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.712 0.000 99.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.712 0.000 99.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.712 0.000 99.864 0.152 ;
    END
  END O1[53]

  PIN O1[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.408 0.000 99.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 99.408 0.000 99.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 99.408 0.000 99.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 99.408 0.000 99.560 0.152 ;
    END
  END O1[52]

  PIN I1[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.192 0.000 98.344 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 98.192 0.000 98.344 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 98.192 0.000 98.344 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 98.192 0.000 98.344 0.152 ;
    END
  END I1[52]

  PIN I1[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.888 0.000 98.040 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.888 0.000 98.040 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.888 0.000 98.040 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.888 0.000 98.040 0.152 ;
    END
  END I1[53]

  PIN I1[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.584 0.000 97.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.584 0.000 97.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.584 0.000 97.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.584 0.000 97.736 0.152 ;
    END
  END I1[54]

  PIN I1[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 97.280 0.000 97.432 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 97.280 0.000 97.432 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 97.280 0.000 97.432 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 97.280 0.000 97.432 0.152 ;
    END
  END I1[55]

  PIN O1[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.064 0.000 96.216 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 96.064 0.000 96.216 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 96.064 0.000 96.216 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 96.064 0.000 96.216 0.152 ;
    END
  END O1[59]

  PIN O1[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.760 0.000 95.912 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.760 0.000 95.912 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.760 0.000 95.912 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.760 0.000 95.912 0.152 ;
    END
  END O1[58]

  PIN O1[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.456 0.000 95.608 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.456 0.000 95.608 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.456 0.000 95.608 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.456 0.000 95.608 0.152 ;
    END
  END O1[57]

  PIN O1[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.152 0.000 95.304 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 95.152 0.000 95.304 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 95.152 0.000 95.304 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 95.152 0.000 95.304 0.152 ;
    END
  END O1[56]

  PIN I1[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.936 0.000 94.088 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.936 0.000 94.088 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.936 0.000 94.088 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.936 0.000 94.088 0.152 ;
    END
  END I1[56]

  PIN I1[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.632 0.000 93.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.632 0.000 93.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.632 0.000 93.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.632 0.000 93.784 0.152 ;
    END
  END I1[57]

  PIN I1[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.328 0.000 93.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.328 0.000 93.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.328 0.000 93.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.328 0.000 93.480 0.152 ;
    END
  END I1[58]

  PIN I1[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 93.024 0.000 93.176 0.152 ;
    END
  END I1[59]

  PIN O1[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.808 0.000 91.960 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 91.808 0.000 91.960 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 91.808 0.000 91.960 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.808 0.000 91.960 0.152 ;
    END
  END O1[63]

  PIN O1[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.504 0.000 91.656 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 91.504 0.000 91.656 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 91.504 0.000 91.656 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.504 0.000 91.656 0.152 ;
    END
  END O1[62]

  PIN O1[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.200 0.000 91.352 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 91.200 0.000 91.352 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 91.200 0.000 91.352 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 91.200 0.000 91.352 0.152 ;
    END
  END O1[61]

  PIN O1[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.896 0.000 91.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 90.896 0.000 91.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 90.896 0.000 91.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 90.896 0.000 91.048 0.152 ;
    END
  END O1[60]

  PIN I1[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.680 0.000 89.832 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.680 0.000 89.832 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.680 0.000 89.832 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.680 0.000 89.832 0.152 ;
    END
  END I1[60]

  PIN I1[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.376 0.000 89.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.376 0.000 89.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.376 0.000 89.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.376 0.000 89.528 0.152 ;
    END
  END I1[61]

  PIN I1[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.072 0.000 89.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 89.072 0.000 89.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 89.072 0.000 89.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 89.072 0.000 89.224 0.152 ;
    END
  END I1[62]

  PIN I1[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 88.768 0.000 88.920 0.152 ;
    END
  END I1[63]

  PIN O1[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.552 0.000 87.704 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.552 0.000 87.704 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.552 0.000 87.704 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.552 0.000 87.704 0.152 ;
    END
  END O1[67]

  PIN O1[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.248 0.000 87.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 87.248 0.000 87.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 87.248 0.000 87.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 87.248 0.000 87.400 0.152 ;
    END
  END O1[66]

  PIN O1[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.944 0.000 87.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.944 0.000 87.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.944 0.000 87.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.944 0.000 87.096 0.152 ;
    END
  END O1[65]

  PIN O1[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 86.640 0.000 86.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 86.640 0.000 86.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 86.640 0.000 86.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 86.640 0.000 86.792 0.152 ;
    END
  END O1[64]

  PIN I1[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.424 0.000 85.576 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.424 0.000 85.576 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.424 0.000 85.576 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.424 0.000 85.576 0.152 ;
    END
  END I1[64]

  PIN I1[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.120 0.000 85.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 85.120 0.000 85.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 85.120 0.000 85.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 85.120 0.000 85.272 0.152 ;
    END
  END I1[65]

  PIN I1[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.816 0.000 84.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.816 0.000 84.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.816 0.000 84.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.816 0.000 84.968 0.152 ;
    END
  END I1[66]

  PIN I1[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 84.512 0.000 84.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 84.512 0.000 84.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 84.512 0.000 84.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 84.512 0.000 84.664 0.152 ;
    END
  END I1[67]

  PIN O1[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.296 0.000 83.448 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 83.296 0.000 83.448 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 83.296 0.000 83.448 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 83.296 0.000 83.448 0.152 ;
    END
  END O1[71]

  PIN O1[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.992 0.000 83.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.992 0.000 83.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.992 0.000 83.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.992 0.000 83.144 0.152 ;
    END
  END O1[70]

  PIN O1[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.688 0.000 82.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.688 0.000 82.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.688 0.000 82.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.688 0.000 82.840 0.152 ;
    END
  END O1[69]

  PIN O1[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 82.384 0.000 82.536 0.152 ;
    END
  END O1[68]

  PIN I1[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 81.168 0.000 81.320 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 81.168 0.000 81.320 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 81.168 0.000 81.320 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 81.168 0.000 81.320 0.152 ;
    END
  END I1[68]

  PIN I1[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.864 0.000 81.016 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.864 0.000 81.016 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.864 0.000 81.016 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.864 0.000 81.016 0.152 ;
    END
  END I1[69]

  PIN I1[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.560 0.000 80.712 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.560 0.000 80.712 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.560 0.000 80.712 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.560 0.000 80.712 0.152 ;
    END
  END I1[70]

  PIN I1[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.256 0.000 80.408 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 80.256 0.000 80.408 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 80.256 0.000 80.408 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 80.256 0.000 80.408 0.152 ;
    END
  END I1[71]

  PIN O1[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.040 0.000 79.192 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 79.040 0.000 79.192 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 79.040 0.000 79.192 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 79.040 0.000 79.192 0.152 ;
    END
  END O1[75]

  PIN O1[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.736 0.000 78.888 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.736 0.000 78.888 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.736 0.000 78.888 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.736 0.000 78.888 0.152 ;
    END
  END O1[74]

  PIN O1[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.432 0.000 78.584 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.432 0.000 78.584 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.432 0.000 78.584 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.432 0.000 78.584 0.152 ;
    END
  END O1[73]

  PIN O1[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.128 0.000 78.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 78.128 0.000 78.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 78.128 0.000 78.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 78.128 0.000 78.280 0.152 ;
    END
  END O1[72]

  PIN I1[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.912 0.000 77.064 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.912 0.000 77.064 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.912 0.000 77.064 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.912 0.000 77.064 0.152 ;
    END
  END I1[72]

  PIN I1[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.608 0.000 76.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.608 0.000 76.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.608 0.000 76.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.608 0.000 76.760 0.152 ;
    END
  END I1[73]

  PIN I1[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.304 0.000 76.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.304 0.000 76.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.304 0.000 76.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.304 0.000 76.456 0.152 ;
    END
  END I1[74]

  PIN I1[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 76.000 0.000 76.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 76.000 0.000 76.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 76.000 0.000 76.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 76.000 0.000 76.152 0.152 ;
    END
  END I1[75]

  PIN O1[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.784 0.000 74.936 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.784 0.000 74.936 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.784 0.000 74.936 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.784 0.000 74.936 0.152 ;
    END
  END O1[79]

  PIN O1[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.480 0.000 74.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.480 0.000 74.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.480 0.000 74.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.480 0.000 74.632 0.152 ;
    END
  END O1[78]

  PIN O1[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.176 0.000 74.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 74.176 0.000 74.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 74.176 0.000 74.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 74.176 0.000 74.328 0.152 ;
    END
  END O1[77]

  PIN O1[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 73.872 0.000 74.024 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 73.872 0.000 74.024 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 73.872 0.000 74.024 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 73.872 0.000 74.024 0.152 ;
    END
  END O1[76]

  PIN I1[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.656 0.000 72.808 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.656 0.000 72.808 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.656 0.000 72.808 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.656 0.000 72.808 0.152 ;
    END
  END I1[76]

  PIN I1[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.352 0.000 72.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.352 0.000 72.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.352 0.000 72.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.352 0.000 72.504 0.152 ;
    END
  END I1[77]

  PIN I1[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.048 0.000 72.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 72.048 0.000 72.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 72.048 0.000 72.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 72.048 0.000 72.200 0.152 ;
    END
  END I1[78]

  PIN I1[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 71.744 0.000 71.896 0.152 ;
    END
  END I1[79]

  PIN O1[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.528 0.000 70.680 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.528 0.000 70.680 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.528 0.000 70.680 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.528 0.000 70.680 0.152 ;
    END
  END O1[83]

  PIN O1[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 70.224 0.000 70.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 70.224 0.000 70.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 70.224 0.000 70.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 70.224 0.000 70.376 0.152 ;
    END
  END O1[82]

  PIN O1[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.920 0.000 70.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.920 0.000 70.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.920 0.000 70.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.920 0.000 70.072 0.152 ;
    END
  END O1[81]

  PIN O1[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.616 0.000 69.768 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 69.616 0.000 69.768 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 69.616 0.000 69.768 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 69.616 0.000 69.768 0.152 ;
    END
  END O1[80]

  PIN I1[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.400 0.000 68.552 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.400 0.000 68.552 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.400 0.000 68.552 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.400 0.000 68.552 0.152 ;
    END
  END I1[80]

  PIN I1[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 68.096 0.000 68.248 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 68.096 0.000 68.248 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 68.096 0.000 68.248 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 68.096 0.000 68.248 0.152 ;
    END
  END I1[81]

  PIN I1[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.792 0.000 67.944 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.792 0.000 67.944 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.792 0.000 67.944 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.792 0.000 67.944 0.152 ;
    END
  END I1[82]

  PIN I1[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.488 0.000 67.640 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 67.488 0.000 67.640 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 67.488 0.000 67.640 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 67.488 0.000 67.640 0.152 ;
    END
  END I1[83]

  PIN O1[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.272 0.000 66.424 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 66.272 0.000 66.424 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 66.272 0.000 66.424 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 66.272 0.000 66.424 0.152 ;
    END
  END O1[87]

  PIN O1[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.968 0.000 66.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.968 0.000 66.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.968 0.000 66.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.968 0.000 66.120 0.152 ;
    END
  END O1[86]

  PIN O1[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.664 0.000 65.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.664 0.000 65.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.664 0.000 65.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.664 0.000 65.816 0.152 ;
    END
  END O1[85]

  PIN O1[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.360 0.000 65.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 65.360 0.000 65.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 65.360 0.000 65.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 65.360 0.000 65.512 0.152 ;
    END
  END O1[84]

  PIN I1[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.144 0.000 64.296 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 64.144 0.000 64.296 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 64.144 0.000 64.296 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 64.144 0.000 64.296 0.152 ;
    END
  END I1[84]

  PIN I1[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.840 0.000 63.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.840 0.000 63.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.840 0.000 63.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.840 0.000 63.992 0.152 ;
    END
  END I1[85]

  PIN I1[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.536 0.000 63.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.536 0.000 63.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.536 0.000 63.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.536 0.000 63.688 0.152 ;
    END
  END I1[86]

  PIN I1[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.232 0.000 63.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 63.232 0.000 63.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 63.232 0.000 63.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 63.232 0.000 63.384 0.152 ;
    END
  END I1[87]

  PIN O1[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 62.016 0.000 62.168 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 62.016 0.000 62.168 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 62.016 0.000 62.168 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 62.016 0.000 62.168 0.152 ;
    END
  END O1[91]

  PIN O1[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.712 0.000 61.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.712 0.000 61.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.712 0.000 61.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.712 0.000 61.864 0.152 ;
    END
  END O1[90]

  PIN O1[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.408 0.000 61.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.408 0.000 61.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.408 0.000 61.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.408 0.000 61.560 0.152 ;
    END
  END O1[89]

  PIN O1[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.104 0.000 61.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 61.104 0.000 61.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 61.104 0.000 61.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 61.104 0.000 61.256 0.152 ;
    END
  END O1[88]

  PIN I1[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.888 0.000 60.040 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.888 0.000 60.040 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.888 0.000 60.040 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.888 0.000 60.040 0.152 ;
    END
  END I1[88]

  PIN I1[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.584 0.000 59.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.584 0.000 59.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.584 0.000 59.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.584 0.000 59.736 0.152 ;
    END
  END I1[89]

  PIN I1[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.280 0.000 59.432 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 59.280 0.000 59.432 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 59.280 0.000 59.432 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 59.280 0.000 59.432 0.152 ;
    END
  END I1[90]

  PIN I1[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.976 0.000 59.128 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 58.976 0.000 59.128 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 58.976 0.000 59.128 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 58.976 0.000 59.128 0.152 ;
    END
  END I1[91]

  PIN O1[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.760 0.000 57.912 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.760 0.000 57.912 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.760 0.000 57.912 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.760 0.000 57.912 0.152 ;
    END
  END O1[95]

  PIN O1[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.456 0.000 57.608 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.456 0.000 57.608 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.456 0.000 57.608 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.456 0.000 57.608 0.152 ;
    END
  END O1[94]

  PIN O1[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.152 0.000 57.304 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 57.152 0.000 57.304 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 57.152 0.000 57.304 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 57.152 0.000 57.304 0.152 ;
    END
  END O1[93]

  PIN O1[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.848 0.000 57.000 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 56.848 0.000 57.000 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 56.848 0.000 57.000 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 56.848 0.000 57.000 0.152 ;
    END
  END O1[92]

  PIN I1[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.632 0.000 55.784 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.632 0.000 55.784 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.632 0.000 55.784 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.632 0.000 55.784 0.152 ;
    END
  END I1[92]

  PIN I1[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.328 0.000 55.480 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.328 0.000 55.480 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.328 0.000 55.480 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.328 0.000 55.480 0.152 ;
    END
  END I1[93]

  PIN I1[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.024 0.000 55.176 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 55.024 0.000 55.176 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 55.024 0.000 55.176 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 55.024 0.000 55.176 0.152 ;
    END
  END I1[94]

  PIN I1[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 54.720 0.000 54.872 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 54.720 0.000 54.872 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 54.720 0.000 54.872 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 54.720 0.000 54.872 0.152 ;
    END
  END I1[95]

  PIN O1[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.504 0.000 53.656 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.504 0.000 53.656 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.504 0.000 53.656 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.504 0.000 53.656 0.152 ;
    END
  END O1[99]

  PIN O1[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.200 0.000 53.352 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 53.200 0.000 53.352 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 53.200 0.000 53.352 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 53.200 0.000 53.352 0.152 ;
    END
  END O1[98]

  PIN O1[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.896 0.000 53.048 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.896 0.000 53.048 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.896 0.000 53.048 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.896 0.000 53.048 0.152 ;
    END
  END O1[97]

  PIN O1[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 52.592 0.000 52.744 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 52.592 0.000 52.744 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 52.592 0.000 52.744 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 52.592 0.000 52.744 0.152 ;
    END
  END O1[96]

  PIN I1[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.376 0.000 51.528 0.152 ;
    END
  END I1[96]

  PIN I1[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 51.072 0.000 51.224 0.152 ;
    END
  END I1[97]

  PIN I1[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.768 0.000 50.920 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.768 0.000 50.920 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.768 0.000 50.920 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.768 0.000 50.920 0.152 ;
    END
  END I1[98]

  PIN I1[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 50.464 0.000 50.616 0.152 ;
    END
  END I1[99]

  PIN O1[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 49.248 0.000 49.400 0.152 ;
    END
  END O1[103]

  PIN O1[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.944 0.000 49.096 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.944 0.000 49.096 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.944 0.000 49.096 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.944 0.000 49.096 0.152 ;
    END
  END O1[102]

  PIN O1[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.640 0.000 48.792 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.640 0.000 48.792 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.640 0.000 48.792 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.640 0.000 48.792 0.152 ;
    END
  END O1[101]

  PIN O1[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.336 0.000 48.488 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 48.336 0.000 48.488 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 48.336 0.000 48.488 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 48.336 0.000 48.488 0.152 ;
    END
  END O1[100]

  PIN I1[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 47.120 0.000 47.272 0.152 ;
    END
  END I1[100]

  PIN I1[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.816 0.000 46.968 0.152 ;
    END
  END I1[101]

  PIN I1[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.512 0.000 46.664 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.512 0.000 46.664 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.512 0.000 46.664 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.512 0.000 46.664 0.152 ;
    END
  END I1[102]

  PIN I1[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 46.208 0.000 46.360 0.152 ;
    END
  END I1[103]

  PIN O1[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.992 0.000 45.144 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.992 0.000 45.144 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.992 0.000 45.144 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.992 0.000 45.144 0.152 ;
    END
  END O1[107]

  PIN O1[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.688 0.000 44.840 0.152 ;
    END
  END O1[106]

  PIN O1[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.384 0.000 44.536 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.384 0.000 44.536 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.384 0.000 44.536 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.384 0.000 44.536 0.152 ;
    END
  END O1[105]

  PIN O1[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 44.080 0.000 44.232 0.152 ;
    END
  END O1[104]

  PIN I1[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.864 0.000 43.016 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.864 0.000 43.016 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.864 0.000 43.016 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.864 0.000 43.016 0.152 ;
    END
  END I1[104]

  PIN I1[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.560 0.000 42.712 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.560 0.000 42.712 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.560 0.000 42.712 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.560 0.000 42.712 0.152 ;
    END
  END I1[105]

  PIN I1[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.256 0.000 42.408 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 42.256 0.000 42.408 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 42.256 0.000 42.408 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 42.256 0.000 42.408 0.152 ;
    END
  END I1[106]

  PIN I1[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.952 0.000 42.104 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 41.952 0.000 42.104 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 41.952 0.000 42.104 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 41.952 0.000 42.104 0.152 ;
    END
  END I1[107]

  PIN O1[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.736 0.000 40.888 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.736 0.000 40.888 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.736 0.000 40.888 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.736 0.000 40.888 0.152 ;
    END
  END O1[111]

  PIN O1[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.432 0.000 40.584 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.432 0.000 40.584 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.432 0.000 40.584 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.432 0.000 40.584 0.152 ;
    END
  END O1[110]

  PIN O1[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.128 0.000 40.280 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 40.128 0.000 40.280 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 40.128 0.000 40.280 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 40.128 0.000 40.280 0.152 ;
    END
  END O1[109]

  PIN O1[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.824 0.000 39.976 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 39.824 0.000 39.976 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 39.824 0.000 39.976 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 39.824 0.000 39.976 0.152 ;
    END
  END O1[108]

  PIN I1[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.608 0.000 38.760 0.152 ;
    END
  END I1[108]

  PIN I1[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.304 0.000 38.456 0.152 ;
    END
  END I1[109]

  PIN I1[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 38.000 0.000 38.152 0.152 ;
    END
  END I1[110]

  PIN I1[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 37.696 0.000 37.848 0.152 ;
    END
  END I1[111]

  PIN O1[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.480 0.000 36.632 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.480 0.000 36.632 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.480 0.000 36.632 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.480 0.000 36.632 0.152 ;
    END
  END O1[115]

  PIN O1[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 36.176 0.000 36.328 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 36.176 0.000 36.328 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 36.176 0.000 36.328 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 36.176 0.000 36.328 0.152 ;
    END
  END O1[114]

  PIN O1[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.872 0.000 36.024 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.872 0.000 36.024 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.872 0.000 36.024 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.872 0.000 36.024 0.152 ;
    END
  END O1[113]

  PIN O1[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.568 0.000 35.720 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 35.568 0.000 35.720 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 35.568 0.000 35.720 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 35.568 0.000 35.720 0.152 ;
    END
  END O1[112]

  PIN I1[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.352 0.000 34.504 0.152 ;
    END
  END I1[112]

  PIN I1[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 34.048 0.000 34.200 0.152 ;
    END
  END I1[113]

  PIN I1[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.744 0.000 33.896 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.744 0.000 33.896 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.744 0.000 33.896 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.744 0.000 33.896 0.152 ;
    END
  END I1[114]

  PIN I1[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.440 0.000 33.592 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 33.440 0.000 33.592 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 33.440 0.000 33.592 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 33.440 0.000 33.592 0.152 ;
    END
  END I1[115]

  PIN O1[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.224 0.000 32.376 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 32.224 0.000 32.376 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 32.224 0.000 32.376 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 32.224 0.000 32.376 0.152 ;
    END
  END O1[119]

  PIN O1[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.920 0.000 32.072 0.152 ;
    END
  END O1[118]

  PIN O1[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.616 0.000 31.768 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.616 0.000 31.768 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.616 0.000 31.768 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.616 0.000 31.768 0.152 ;
    END
  END O1[117]

  PIN O1[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.312 0.000 31.464 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 31.312 0.000 31.464 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 31.312 0.000 31.464 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 31.312 0.000 31.464 0.152 ;
    END
  END O1[116]

  PIN I1[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 30.096 0.000 30.248 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 30.096 0.000 30.248 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 30.096 0.000 30.248 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 30.096 0.000 30.248 0.152 ;
    END
  END I1[116]

  PIN I1[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.792 0.000 29.944 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.792 0.000 29.944 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.792 0.000 29.944 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.792 0.000 29.944 0.152 ;
    END
  END I1[117]

  PIN I1[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.488 0.000 29.640 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.488 0.000 29.640 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.488 0.000 29.640 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.488 0.000 29.640 0.152 ;
    END
  END I1[118]

  PIN I1[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.184 0.000 29.336 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 29.184 0.000 29.336 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 29.184 0.000 29.336 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 29.184 0.000 29.336 0.152 ;
    END
  END I1[119]

  PIN O1[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.968 0.000 28.120 0.152 ;
    END
  END O1[123]

  PIN O1[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.664 0.000 27.816 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.664 0.000 27.816 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.664 0.000 27.816 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.664 0.000 27.816 0.152 ;
    END
  END O1[122]

  PIN O1[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.360 0.000 27.512 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.360 0.000 27.512 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.360 0.000 27.512 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.360 0.000 27.512 0.152 ;
    END
  END O1[121]

  PIN O1[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.056 0.000 27.208 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 27.056 0.000 27.208 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 27.056 0.000 27.208 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 27.056 0.000 27.208 0.152 ;
    END
  END O1[120]

  PIN I1[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.840 0.000 25.992 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.840 0.000 25.992 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.840 0.000 25.992 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.840 0.000 25.992 0.152 ;
    END
  END I1[120]

  PIN I1[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.536 0.000 25.688 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.536 0.000 25.688 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.536 0.000 25.688 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.536 0.000 25.688 0.152 ;
    END
  END I1[121]

  PIN I1[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 25.232 0.000 25.384 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 25.232 0.000 25.384 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 25.232 0.000 25.384 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 25.232 0.000 25.384 0.152 ;
    END
  END I1[122]

  PIN I1[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.928 0.000 25.080 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 24.928 0.000 25.080 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 24.928 0.000 25.080 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 24.928 0.000 25.080 0.152 ;
    END
  END I1[123]

  PIN O1[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.712 0.000 23.864 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.712 0.000 23.864 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.712 0.000 23.864 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.712 0.000 23.864 0.152 ;
    END
  END O1[127]

  PIN O1[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.408 0.000 23.560 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.408 0.000 23.560 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.408 0.000 23.560 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.408 0.000 23.560 0.152 ;
    END
  END O1[126]

  PIN O1[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.104 0.000 23.256 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 23.104 0.000 23.256 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 23.104 0.000 23.256 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 23.104 0.000 23.256 0.152 ;
    END
  END O1[125]

  PIN O1[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.800 0.000 22.952 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 22.800 0.000 22.952 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 22.800 0.000 22.952 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 22.800 0.000 22.952 0.152 ;
    END
  END O1[124]

  PIN I1[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.584 0.000 21.736 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.584 0.000 21.736 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.584 0.000 21.736 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.584 0.000 21.736 0.152 ;
    END
  END I1[124]

  PIN I1[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.280 0.000 21.432 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 21.280 0.000 21.432 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 21.280 0.000 21.432 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 21.280 0.000 21.432 0.152 ;
    END
  END I1[125]

  PIN I1[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.976 0.000 21.128 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.976 0.000 21.128 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.976 0.000 21.128 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.976 0.000 21.128 0.152 ;
    END
  END I1[126]

  PIN I1[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 20.672 0.000 20.824 0.152 ;
    END
    PORT
      LAYER M3 ;
        RECT 20.672 0.000 20.824 0.152 ;
    END
    PORT
      LAYER M4 ;
        RECT 20.672 0.000 20.824 0.152 ;
    END
    PORT
      LAYER M5 ;
        RECT 20.672 0.000 20.824 0.152 ;
    END
  END I1[127]

  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.384 85.120 177.536 85.272 ;
    END
    PORT
      LAYER M3 ;
        RECT 177.384 85.120 177.536 85.272 ;
    END
    PORT
      LAYER M4 ;
        RECT 177.384 85.120 177.536 85.272 ;
    END
    PORT
      LAYER M5 ;
        RECT 177.384 85.120 177.536 85.272 ;
    END
  END A1[0]

  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.384 81.472 177.536 81.624 ;
    END
    PORT
      LAYER M3 ;
        RECT 177.384 81.472 177.536 81.624 ;
    END
    PORT
      LAYER M4 ;
        RECT 177.384 81.472 177.536 81.624 ;
    END
    PORT
      LAYER M5 ;
        RECT 177.384 81.472 177.536 81.624 ;
    END
  END A1[1]

  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.384 77.824 177.536 77.976 ;
    END
    PORT
      LAYER M3 ;
        RECT 177.384 77.824 177.536 77.976 ;
    END
    PORT
      LAYER M4 ;
        RECT 177.384 77.824 177.536 77.976 ;
    END
    PORT
      LAYER M5 ;
        RECT 177.384 77.824 177.536 77.976 ;
    END
  END A1[2]

  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.384 74.176 177.536 74.328 ;
    END
    PORT
      LAYER M3 ;
        RECT 177.384 74.176 177.536 74.328 ;
    END
    PORT
      LAYER M4 ;
        RECT 177.384 74.176 177.536 74.328 ;
    END
    PORT
      LAYER M5 ;
        RECT 177.384 74.176 177.536 74.328 ;
    END
  END A1[3]

  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.384 70.528 177.536 70.680 ;
    END
    PORT
      LAYER M3 ;
        RECT 177.384 70.528 177.536 70.680 ;
    END
    PORT
      LAYER M4 ;
        RECT 177.384 70.528 177.536 70.680 ;
    END
    PORT
      LAYER M5 ;
        RECT 177.384 70.528 177.536 70.680 ;
    END
  END A1[4]

  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.384 66.880 177.536 67.032 ;
    END
    PORT
      LAYER M3 ;
        RECT 177.384 66.880 177.536 67.032 ;
    END
    PORT
      LAYER M4 ;
        RECT 177.384 66.880 177.536 67.032 ;
    END
    PORT
      LAYER M5 ;
        RECT 177.384 66.880 177.536 67.032 ;
    END
  END A1[5]

  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.384 63.232 177.536 63.384 ;
    END
    PORT
      LAYER M3 ;
        RECT 177.384 63.232 177.536 63.384 ;
    END
    PORT
      LAYER M4 ;
        RECT 177.384 63.232 177.536 63.384 ;
    END
    PORT
      LAYER M5 ;
        RECT 177.384 63.232 177.536 63.384 ;
    END
  END A1[6]

  PIN A1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.384 59.584 177.536 59.736 ;
    END
    PORT
      LAYER M3 ;
        RECT 177.384 59.584 177.536 59.736 ;
    END
    PORT
      LAYER M4 ;
        RECT 177.384 59.584 177.536 59.736 ;
    END
    PORT
      LAYER M5 ;
        RECT 177.384 59.584 177.536 59.736 ;
    END
  END A1[7]

  PIN A1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.384 55.936 177.536 56.088 ;
    END
    PORT
      LAYER M3 ;
        RECT 177.384 55.936 177.536 56.088 ;
    END
    PORT
      LAYER M4 ;
        RECT 177.384 55.936 177.536 56.088 ;
    END
    PORT
      LAYER M5 ;
        RECT 177.384 55.936 177.536 56.088 ;
    END
  END A1[8]

  PIN WEB1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 177.384 24.320 177.536 24.472 ;
    END
    PORT
      LAYER M3 ;
        RECT 177.384 24.320 177.536 24.472 ;
    END
    PORT
      LAYER M4 ;
        RECT 177.384 24.320 177.536 24.472 ;
    END
    PORT
      LAYER M5 ;
        RECT 177.384 24.320 177.536 24.472 ;
    END
  END WEB1

  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M2 ;
        RECT 5.195 95.280 7.195 97.280 ;
    END
    PORT
      LAYER M3 ;
        RECT 5.195 95.280 7.195 97.280 ;
    END
    PORT
      LAYER M5 ;
        RECT 5.195 95.280 7.195 97.280 ;
    END
  END VDD

  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M2 ;
        RECT 7.915 95.280 9.915 97.280 ;
    END
    PORT
      LAYER M3 ;
        RECT 7.915 95.280 9.915 97.280 ;
    END
    PORT
      LAYER M5 ;
        RECT 7.915 95.280 9.915 97.280 ;
    END
  END VSS

  OBS
    LAYER M2 ;
      RECT 159.600 0.000 177.536 0.304 ;
      RECT 158.384 0.000 159.144 0.304 ;
      RECT 157.168 0.000 157.928 0.304 ;
      RECT 155.952 0.000 156.712 0.304 ;
      RECT 153.824 0.000 154.584 0.304 ;
      RECT 151.696 0.000 152.456 0.304 ;
      RECT 149.568 0.000 150.328 0.304 ;
      RECT 147.440 0.000 148.200 0.304 ;
      RECT 145.312 0.000 146.072 0.304 ;
      RECT 143.184 0.000 143.944 0.304 ;
      RECT 141.056 0.000 141.816 0.304 ;
      RECT 138.928 0.000 139.688 0.304 ;
      RECT 136.800 0.000 137.560 0.304 ;
      RECT 134.672 0.000 135.432 0.304 ;
      RECT 132.544 0.000 133.304 0.304 ;
      RECT 130.416 0.000 131.176 0.304 ;
      RECT 128.288 0.000 129.048 0.304 ;
      RECT 126.160 0.000 126.920 0.304 ;
      RECT 124.032 0.000 124.792 0.304 ;
      RECT 121.904 0.000 122.664 0.304 ;
      RECT 119.776 0.000 120.536 0.304 ;
      RECT 117.648 0.000 118.408 0.304 ;
      RECT 115.520 0.000 116.280 0.304 ;
      RECT 113.392 0.000 114.152 0.304 ;
      RECT 111.264 0.000 112.024 0.304 ;
      RECT 109.136 0.000 109.896 0.304 ;
      RECT 107.008 0.000 107.768 0.304 ;
      RECT 104.880 0.000 105.640 0.304 ;
      RECT 102.752 0.000 103.512 0.304 ;
      RECT 100.624 0.000 101.384 0.304 ;
      RECT 98.496 0.000 99.256 0.304 ;
      RECT 96.368 0.000 97.128 0.304 ;
      RECT 94.240 0.000 95.000 0.304 ;
      RECT 92.112 0.000 92.872 0.304 ;
      RECT 89.984 0.000 90.744 0.304 ;
      RECT 87.856 0.000 88.616 0.304 ;
      RECT 85.728 0.000 86.488 0.304 ;
      RECT 83.600 0.000 84.360 0.304 ;
      RECT 81.472 0.000 82.232 0.304 ;
      RECT 79.344 0.000 80.104 0.304 ;
      RECT 77.216 0.000 77.976 0.304 ;
      RECT 75.088 0.000 75.848 0.304 ;
      RECT 72.960 0.000 73.720 0.304 ;
      RECT 70.832 0.000 71.592 0.304 ;
      RECT 68.704 0.000 69.464 0.304 ;
      RECT 66.576 0.000 67.336 0.304 ;
      RECT 64.448 0.000 65.208 0.304 ;
      RECT 62.320 0.000 63.080 0.304 ;
      RECT 60.192 0.000 60.952 0.304 ;
      RECT 58.064 0.000 58.824 0.304 ;
      RECT 55.936 0.000 56.696 0.304 ;
      RECT 53.808 0.000 54.568 0.304 ;
      RECT 51.680 0.000 52.440 0.304 ;
      RECT 49.552 0.000 50.312 0.304 ;
      RECT 47.424 0.000 48.184 0.304 ;
      RECT 45.296 0.000 46.056 0.304 ;
      RECT 43.168 0.000 43.928 0.304 ;
      RECT 41.040 0.000 41.800 0.304 ;
      RECT 38.912 0.000 39.672 0.304 ;
      RECT 36.784 0.000 37.544 0.304 ;
      RECT 34.656 0.000 35.416 0.304 ;
      RECT 32.528 0.000 33.288 0.304 ;
      RECT 30.400 0.000 31.160 0.304 ;
      RECT 28.272 0.000 29.032 0.304 ;
      RECT 26.144 0.000 26.904 0.304 ;
      RECT 24.016 0.000 24.776 0.304 ;
      RECT 21.888 0.000 22.648 0.304 ;
      RECT 0.000 0.000 20.520 0.304 ;
      RECT 177.232 85.424 177.536 95.128 ;
      RECT 177.232 81.776 177.536 84.968 ;
      RECT 177.232 78.128 177.536 81.320 ;
      RECT 177.232 74.480 177.536 77.672 ;
      RECT 177.232 70.832 177.536 74.024 ;
      RECT 177.232 67.184 177.536 70.376 ;
      RECT 177.232 63.536 177.536 66.728 ;
      RECT 177.232 59.888 177.536 63.080 ;
      RECT 177.232 56.240 177.536 59.432 ;
      RECT 177.232 24.624 177.536 55.784 ;
      RECT 177.232 0.304 177.536 24.168 ;
      RECT 0.000 95.128 5.043 97.280 ;
      RECT 7.355 95.128 7.763 97.280 ;
      RECT 10.067 95.128 177.536 97.280 ;
      RECT 0.000 0.304 177.232 95.128 ;
    LAYER M3 ;
      RECT 159.600 0.000 177.536 0.304 ;
      RECT 158.384 0.000 159.144 0.304 ;
      RECT 157.168 0.000 157.928 0.304 ;
      RECT 155.952 0.000 156.712 0.304 ;
      RECT 153.824 0.000 154.584 0.304 ;
      RECT 151.696 0.000 152.456 0.304 ;
      RECT 149.568 0.000 150.328 0.304 ;
      RECT 147.440 0.000 148.200 0.304 ;
      RECT 145.312 0.000 146.072 0.304 ;
      RECT 143.184 0.000 143.944 0.304 ;
      RECT 141.056 0.000 141.816 0.304 ;
      RECT 138.928 0.000 139.688 0.304 ;
      RECT 136.800 0.000 137.560 0.304 ;
      RECT 134.672 0.000 135.432 0.304 ;
      RECT 132.544 0.000 133.304 0.304 ;
      RECT 130.416 0.000 131.176 0.304 ;
      RECT 128.288 0.000 129.048 0.304 ;
      RECT 126.160 0.000 126.920 0.304 ;
      RECT 124.032 0.000 124.792 0.304 ;
      RECT 121.904 0.000 122.664 0.304 ;
      RECT 119.776 0.000 120.536 0.304 ;
      RECT 117.648 0.000 118.408 0.304 ;
      RECT 115.520 0.000 116.280 0.304 ;
      RECT 113.392 0.000 114.152 0.304 ;
      RECT 111.264 0.000 112.024 0.304 ;
      RECT 109.136 0.000 109.896 0.304 ;
      RECT 107.008 0.000 107.768 0.304 ;
      RECT 104.880 0.000 105.640 0.304 ;
      RECT 102.752 0.000 103.512 0.304 ;
      RECT 100.624 0.000 101.384 0.304 ;
      RECT 98.496 0.000 99.256 0.304 ;
      RECT 96.368 0.000 97.128 0.304 ;
      RECT 94.240 0.000 95.000 0.304 ;
      RECT 92.112 0.000 92.872 0.304 ;
      RECT 89.984 0.000 90.744 0.304 ;
      RECT 87.856 0.000 88.616 0.304 ;
      RECT 85.728 0.000 86.488 0.304 ;
      RECT 83.600 0.000 84.360 0.304 ;
      RECT 81.472 0.000 82.232 0.304 ;
      RECT 79.344 0.000 80.104 0.304 ;
      RECT 77.216 0.000 77.976 0.304 ;
      RECT 75.088 0.000 75.848 0.304 ;
      RECT 72.960 0.000 73.720 0.304 ;
      RECT 70.832 0.000 71.592 0.304 ;
      RECT 68.704 0.000 69.464 0.304 ;
      RECT 66.576 0.000 67.336 0.304 ;
      RECT 64.448 0.000 65.208 0.304 ;
      RECT 62.320 0.000 63.080 0.304 ;
      RECT 60.192 0.000 60.952 0.304 ;
      RECT 58.064 0.000 58.824 0.304 ;
      RECT 55.936 0.000 56.696 0.304 ;
      RECT 53.808 0.000 54.568 0.304 ;
      RECT 51.680 0.000 52.440 0.304 ;
      RECT 49.552 0.000 50.312 0.304 ;
      RECT 47.424 0.000 48.184 0.304 ;
      RECT 45.296 0.000 46.056 0.304 ;
      RECT 43.168 0.000 43.928 0.304 ;
      RECT 41.040 0.000 41.800 0.304 ;
      RECT 38.912 0.000 39.672 0.304 ;
      RECT 36.784 0.000 37.544 0.304 ;
      RECT 34.656 0.000 35.416 0.304 ;
      RECT 32.528 0.000 33.288 0.304 ;
      RECT 30.400 0.000 31.160 0.304 ;
      RECT 28.272 0.000 29.032 0.304 ;
      RECT 26.144 0.000 26.904 0.304 ;
      RECT 24.016 0.000 24.776 0.304 ;
      RECT 21.888 0.000 22.648 0.304 ;
      RECT 0.000 0.000 20.520 0.304 ;
      RECT 177.232 85.424 177.536 95.128 ;
      RECT 177.232 81.776 177.536 84.968 ;
      RECT 177.232 78.128 177.536 81.320 ;
      RECT 177.232 74.480 177.536 77.672 ;
      RECT 177.232 70.832 177.536 74.024 ;
      RECT 177.232 67.184 177.536 70.376 ;
      RECT 177.232 63.536 177.536 66.728 ;
      RECT 177.232 59.888 177.536 63.080 ;
      RECT 177.232 56.240 177.536 59.432 ;
      RECT 177.232 24.624 177.536 55.784 ;
      RECT 177.232 0.304 177.536 24.168 ;
      RECT 0.000 95.128 5.043 97.280 ;
      RECT 7.355 95.128 7.763 97.280 ;
      RECT 10.067 95.128 177.536 97.280 ;
      RECT 0.000 0.304 177.232 95.128 ;
    LAYER M4 ;
      RECT 159.600 0.000 177.536 0.304 ;
      RECT 158.384 0.000 159.144 0.304 ;
      RECT 157.168 0.000 157.928 0.304 ;
      RECT 155.952 0.000 156.712 0.304 ;
      RECT 153.824 0.000 154.584 0.304 ;
      RECT 151.696 0.000 152.456 0.304 ;
      RECT 149.568 0.000 150.328 0.304 ;
      RECT 147.440 0.000 148.200 0.304 ;
      RECT 145.312 0.000 146.072 0.304 ;
      RECT 143.184 0.000 143.944 0.304 ;
      RECT 141.056 0.000 141.816 0.304 ;
      RECT 138.928 0.000 139.688 0.304 ;
      RECT 136.800 0.000 137.560 0.304 ;
      RECT 134.672 0.000 135.432 0.304 ;
      RECT 132.544 0.000 133.304 0.304 ;
      RECT 130.416 0.000 131.176 0.304 ;
      RECT 128.288 0.000 129.048 0.304 ;
      RECT 126.160 0.000 126.920 0.304 ;
      RECT 124.032 0.000 124.792 0.304 ;
      RECT 121.904 0.000 122.664 0.304 ;
      RECT 119.776 0.000 120.536 0.304 ;
      RECT 117.648 0.000 118.408 0.304 ;
      RECT 115.520 0.000 116.280 0.304 ;
      RECT 113.392 0.000 114.152 0.304 ;
      RECT 111.264 0.000 112.024 0.304 ;
      RECT 109.136 0.000 109.896 0.304 ;
      RECT 107.008 0.000 107.768 0.304 ;
      RECT 104.880 0.000 105.640 0.304 ;
      RECT 102.752 0.000 103.512 0.304 ;
      RECT 100.624 0.000 101.384 0.304 ;
      RECT 98.496 0.000 99.256 0.304 ;
      RECT 96.368 0.000 97.128 0.304 ;
      RECT 94.240 0.000 95.000 0.304 ;
      RECT 92.112 0.000 92.872 0.304 ;
      RECT 89.984 0.000 90.744 0.304 ;
      RECT 87.856 0.000 88.616 0.304 ;
      RECT 85.728 0.000 86.488 0.304 ;
      RECT 83.600 0.000 84.360 0.304 ;
      RECT 81.472 0.000 82.232 0.304 ;
      RECT 79.344 0.000 80.104 0.304 ;
      RECT 77.216 0.000 77.976 0.304 ;
      RECT 75.088 0.000 75.848 0.304 ;
      RECT 72.960 0.000 73.720 0.304 ;
      RECT 70.832 0.000 71.592 0.304 ;
      RECT 68.704 0.000 69.464 0.304 ;
      RECT 66.576 0.000 67.336 0.304 ;
      RECT 64.448 0.000 65.208 0.304 ;
      RECT 62.320 0.000 63.080 0.304 ;
      RECT 60.192 0.000 60.952 0.304 ;
      RECT 58.064 0.000 58.824 0.304 ;
      RECT 55.936 0.000 56.696 0.304 ;
      RECT 53.808 0.000 54.568 0.304 ;
      RECT 51.680 0.000 52.440 0.304 ;
      RECT 49.552 0.000 50.312 0.304 ;
      RECT 47.424 0.000 48.184 0.304 ;
      RECT 45.296 0.000 46.056 0.304 ;
      RECT 43.168 0.000 43.928 0.304 ;
      RECT 41.040 0.000 41.800 0.304 ;
      RECT 38.912 0.000 39.672 0.304 ;
      RECT 36.784 0.000 37.544 0.304 ;
      RECT 34.656 0.000 35.416 0.304 ;
      RECT 32.528 0.000 33.288 0.304 ;
      RECT 30.400 0.000 31.160 0.304 ;
      RECT 28.272 0.000 29.032 0.304 ;
      RECT 26.144 0.000 26.904 0.304 ;
      RECT 24.016 0.000 24.776 0.304 ;
      RECT 21.888 0.000 22.648 0.304 ;
      RECT 0.000 0.000 20.520 0.304 ;
      RECT 177.232 85.424 177.536 95.128 ;
      RECT 177.232 81.776 177.536 84.968 ;
      RECT 177.232 78.128 177.536 81.320 ;
      RECT 177.232 74.480 177.536 77.672 ;
      RECT 177.232 70.832 177.536 74.024 ;
      RECT 177.232 67.184 177.536 70.376 ;
      RECT 177.232 63.536 177.536 66.728 ;
      RECT 177.232 59.888 177.536 63.080 ;
      RECT 177.232 56.240 177.536 59.432 ;
      RECT 177.232 24.624 177.536 55.784 ;
      RECT 177.232 0.304 177.536 24.168 ;
      RECT 0.000 95.128 5.043 97.280 ;
      RECT 7.355 95.128 7.763 97.280 ;
      RECT 10.067 95.128 177.536 97.280 ;
      RECT 0.000 0.304 177.232 95.128 ;
    LAYER M5 ;
      RECT 159.600 0.000 177.536 0.304 ;
      RECT 158.384 0.000 159.144 0.304 ;
      RECT 157.168 0.000 157.928 0.304 ;
      RECT 155.952 0.000 156.712 0.304 ;
      RECT 153.824 0.000 154.584 0.304 ;
      RECT 151.696 0.000 152.456 0.304 ;
      RECT 149.568 0.000 150.328 0.304 ;
      RECT 147.440 0.000 148.200 0.304 ;
      RECT 145.312 0.000 146.072 0.304 ;
      RECT 143.184 0.000 143.944 0.304 ;
      RECT 141.056 0.000 141.816 0.304 ;
      RECT 138.928 0.000 139.688 0.304 ;
      RECT 136.800 0.000 137.560 0.304 ;
      RECT 134.672 0.000 135.432 0.304 ;
      RECT 132.544 0.000 133.304 0.304 ;
      RECT 130.416 0.000 131.176 0.304 ;
      RECT 128.288 0.000 129.048 0.304 ;
      RECT 126.160 0.000 126.920 0.304 ;
      RECT 124.032 0.000 124.792 0.304 ;
      RECT 121.904 0.000 122.664 0.304 ;
      RECT 119.776 0.000 120.536 0.304 ;
      RECT 117.648 0.000 118.408 0.304 ;
      RECT 115.520 0.000 116.280 0.304 ;
      RECT 113.392 0.000 114.152 0.304 ;
      RECT 111.264 0.000 112.024 0.304 ;
      RECT 109.136 0.000 109.896 0.304 ;
      RECT 107.008 0.000 107.768 0.304 ;
      RECT 104.880 0.000 105.640 0.304 ;
      RECT 102.752 0.000 103.512 0.304 ;
      RECT 100.624 0.000 101.384 0.304 ;
      RECT 98.496 0.000 99.256 0.304 ;
      RECT 96.368 0.000 97.128 0.304 ;
      RECT 94.240 0.000 95.000 0.304 ;
      RECT 92.112 0.000 92.872 0.304 ;
      RECT 89.984 0.000 90.744 0.304 ;
      RECT 87.856 0.000 88.616 0.304 ;
      RECT 85.728 0.000 86.488 0.304 ;
      RECT 83.600 0.000 84.360 0.304 ;
      RECT 81.472 0.000 82.232 0.304 ;
      RECT 79.344 0.000 80.104 0.304 ;
      RECT 77.216 0.000 77.976 0.304 ;
      RECT 75.088 0.000 75.848 0.304 ;
      RECT 72.960 0.000 73.720 0.304 ;
      RECT 70.832 0.000 71.592 0.304 ;
      RECT 68.704 0.000 69.464 0.304 ;
      RECT 66.576 0.000 67.336 0.304 ;
      RECT 64.448 0.000 65.208 0.304 ;
      RECT 62.320 0.000 63.080 0.304 ;
      RECT 60.192 0.000 60.952 0.304 ;
      RECT 58.064 0.000 58.824 0.304 ;
      RECT 55.936 0.000 56.696 0.304 ;
      RECT 53.808 0.000 54.568 0.304 ;
      RECT 51.680 0.000 52.440 0.304 ;
      RECT 49.552 0.000 50.312 0.304 ;
      RECT 47.424 0.000 48.184 0.304 ;
      RECT 45.296 0.000 46.056 0.304 ;
      RECT 43.168 0.000 43.928 0.304 ;
      RECT 41.040 0.000 41.800 0.304 ;
      RECT 38.912 0.000 39.672 0.304 ;
      RECT 36.784 0.000 37.544 0.304 ;
      RECT 34.656 0.000 35.416 0.304 ;
      RECT 32.528 0.000 33.288 0.304 ;
      RECT 30.400 0.000 31.160 0.304 ;
      RECT 28.272 0.000 29.032 0.304 ;
      RECT 26.144 0.000 26.904 0.304 ;
      RECT 24.016 0.000 24.776 0.304 ;
      RECT 21.888 0.000 22.648 0.304 ;
      RECT 0.000 0.000 20.520 0.304 ;
      RECT 177.232 85.424 177.536 95.128 ;
      RECT 177.232 81.776 177.536 84.968 ;
      RECT 177.232 78.128 177.536 81.320 ;
      RECT 177.232 74.480 177.536 77.672 ;
      RECT 177.232 70.832 177.536 74.024 ;
      RECT 177.232 67.184 177.536 70.376 ;
      RECT 177.232 63.536 177.536 66.728 ;
      RECT 177.232 59.888 177.536 63.080 ;
      RECT 177.232 56.240 177.536 59.432 ;
      RECT 177.232 24.624 177.536 55.784 ;
      RECT 177.232 0.304 177.536 24.168 ;
      RECT 0.000 95.128 5.043 97.280 ;
      RECT 7.355 95.128 7.763 97.280 ;
      RECT 10.067 95.128 177.536 97.280 ;
      RECT 0.000 0.304 177.232 95.128 ;
  END

END sram6t512x128

END LIBRARY
